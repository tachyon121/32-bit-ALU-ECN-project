`timescale 1 ns/1 ps
    `include "alu.v"


    module sub_tb ();
        reg clock;
        reg [31:0] x1, x2;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] x3;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .x1(x1),
                .x2(x2),
                .OpCode(op),
                .x3(x3)
            );
        /* create x1 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, x1, x2, op, x3);
            clock = 0;

    op = 3'b001;

		/* Display the operation */
		$display ("Opcode: 001, Operation: SUB");
		/* Test Cases!*/
		x1 = 32'b11111101110101110011001010100000;
		x2 = 32'b01000001010111010111101010010001;
		correct = 32'b11111101110101110011001010100000;
		#400; //-3.575586e+37 * 13.842423 = -3.575586e+37
				
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110011110110110011000101110111;
		x2 = 32'b00011110110111101110001001110110;
		correct = 32'b10110011110110110011000101110111;
		#400; //-1.020698e-07 * 2.3598826e-20 = -1.020698e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100100000001111011110101110;
		x2 = 32'b01011101101110001111011100011101;
		correct = 32'b11011101101110001111011100011101;
		#400; //-3.6654768e-12 * 1.6660192e+18 = -1.6660192e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001101100001110010001010101110;
		x2 = 32'b10110000100000110101110000100100;
		correct = 32'b11001101100001110010001010101110;
		#400; //-283399600.0 * -9.557692e-10 = -283399600.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101110011100110110101101100;
		x2 = 32'b00001101100100110001001011001100;
		correct = 32'b11111101110011100110110101101100;
		#400; //-3.429864e+37 * 9.0641e-31 = -3.429864e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011010010100110010100101010000;
		x2 = 32'b10001110111100100110010111011101;
		correct = 32'b10011010010100110010100101001110;
		#400; //-4.366715e-23 * -5.9755697e-30 = -4.3667143e-23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011010100111011101000101000;
		x2 = 32'b11011110110101101011010101010011;
		correct = 32'b01011110110101101011010101010011;
		#400; //1.1477753e-17 * -7.7356817e+18 = 7.7356817e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001011010111000011101111001;
		x2 = 32'b01011111110110110110000000111111;
		correct = 32'b01111001011010111000011101111001;
		#400; //7.643359e+34 * 3.1615408e+19 = 7.643359e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000001111000001001101110010;
		x2 = 32'b01100111001101110011011011010111;
		correct = 32'b11100111001101110011011011010111;
		#400; //12621564000.0 * 8.652047e+23 = -8.652047e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110100100101110001000011110;
		x2 = 32'b11000101110110011000110101011000;
		correct = 32'b01000101110110011000111110100100;
		#400; //0.2868814 * -6961.668 = 6961.955
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011001010001101110011011100001;
		x2 = 32'b11001011000010011101010011000001;
		correct = 32'b11011001010001101110011011100001;
		#400; //-3499118700000000.0 * -9032897.0 = -3499118700000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011010000000000011010100110;
		x2 = 32'b10101101111010100111011011001011;
		correct = 32'b00101101111010100111011011010001;
		#400; //1.0409749e-17 * -2.6655475e-11 = 2.6655485e-11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101001011011000111100100010101;
		x2 = 32'b11100100100101010000000000110100;
		correct = 32'b11101001011011000010111010010101;
		#400; //-1.7867393e+25 * -2.1988636e+22 = -1.7845404e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011100111010001101010001011101;
		x2 = 32'b11101010100000111000010010111111;
		correct = 32'b01101010100000111000010010111111;
		#400; //-5.2428552e+17 * -7.949808e+25 = 7.949808e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100010000010010101000100110111;
		x2 = 32'b10101101011001111001000101000111;
		correct = 32'b01100010000010010101000100110111;
		#400; //6.33264e+20 * -1.3163088e-11 = 6.33264e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100001111101000011111010110;
		x2 = 32'b01110101001100001110010001001011;
		correct = 32'b11110101000000010100001001010110;
		#400; //6.038156e+31 * 2.2423696e+32 = -1.638554e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100010111011100110000111111111;
		x2 = 32'b01011011110010110011100001101111;
		correct = 32'b11011011110010110011100001101111;
		#400; //6.4613787e-18 * 1.1440294e+17 = -1.1440294e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001110010001001010000100110110;
		x2 = 32'b00001100010110011000000010110000;
		correct = 32'b01001110010001001010000100110110;
		#400; //824724860.0 * 1.6755797e-31 = 824724860.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001001110001111010110001010111;
		x2 = 32'b01100111110111011011101011110011;
		correct = 32'b11100111110111011011101011110011;
		#400; //4.8069575e-33 * 2.0941832e+24 = -2.0941832e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111000110101100001001100100000;
		x2 = 32'b00000111011111101011001110010010;
		correct = 32'b10111000110101100001001100100000;
		#400; //-0.000102078775 * 1.9161607e-34 = -0.000102078775
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100110001110100100110101111000;
		x2 = 32'b10100000000011000110101001010101;
		correct = 32'b11100110001110100100110101111000;
		#400; //-2.199473e+23 * -1.1893644e-19 = -2.199473e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100101101000000100110010001;
		x2 = 32'b01011100000110100000011101111010;
		correct = 32'b11011100000110100000011101111010;
		#400; //-1.8179129e-26 * 1.7342147e+17 = -1.7342147e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110001111000011010010100111;
		x2 = 32'b00011010100101111001111101000010;
		correct = 32'b10011010100101111001111101000010;
		#400; //3.5397553e-35 * 6.270943e-23 = -6.270943e-23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010010000010011011001100110001;
		x2 = 32'b11010001000001000111100000110011;
		correct = 32'b01010001000001000111100000110011;
		#400; //-4.345045e-28 * -35559520000.0 = 35559520000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010101100111100100111110111101;
		x2 = 32'b01110111110101010000111010101101;
		correct = 32'b11110111110101010000111010101101;
		#400; //6.3941497e-26 * 8.642632e+33 = -8.642632e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111100011000001001001001101;
		x2 = 32'b10100010100011000110001000111001;
		correct = 32'b11010111100011000001001001001101;
		#400; //-308020460000000.0 * -3.8051073e-18 = -308020460000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011000010110000110000000010110;
		x2 = 32'b11011011111011001110010101111011;
		correct = 32'b01011011111010110011010010111011;
		#400; //-951628800000000.0 * -1.3336082e+17 = 1.32409195e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011111010100001010000001100101;
		x2 = 32'b01000111001000100010011001111110;
		correct = 32'b11000111001000100010011001111110;
		#400; //-4.417839e-20 * 41510.492 = -41510.492
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101101010001110110011010111110;
		x2 = 32'b01001111001101000110111001100101;
		correct = 32'b11101101010001110110011010111110;
		#400; //-3.8569828e+27 * 3027133700.0 = -3.8569828e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100110110101110111111100101111;
		x2 = 32'b11000001100001010110110101111001;
		correct = 32'b01000001100001010110110101111001;
		#400; //-1.4953095e-15 * -16.678453 = 16.678453
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010011110101100100010101001010;
		x2 = 32'b10101111110110101000010111010111;
		correct = 32'b01010011110101100100010101001010;
		#400; //1840571000000.0 * -3.9749068e-10 = 1840571000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000111111000011010010001101111;
		x2 = 32'b11111111110111001101101100111011;
		correct = 32'b11111111110111001101101100111011;
		#400; //-3.3950883e-34 * nan = nan
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111000101011001110010011001;
		x2 = 32'b00000001011001010111100000011000;
		correct = 32'b10111111000101011001110010011001;
		#400; //-0.58442074 * 4.214682e-38 = -0.58442074
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110101001001101011100000101010;
		x2 = 32'b01101011011110011001001000010100;
		correct = 32'b11101011011110011001001000010100;
		#400; //-6.2107813e-07 * 3.0171236e+26 = -3.0171236e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011110110011001000111110001000;
		x2 = 32'b11110011001101111101001111010110;
		correct = 32'b01110011001101111101001111010110;
		#400; //2.1658703e-20 * -1.4564314e+31 = 1.4564314e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110101111111111001101000001111;
		x2 = 32'b00001011111010011111101101010110;
		correct = 32'b11110101111111111001101000001111;
		#400; //-6.4802753e+32 * 9.0126504e-32 = -6.4802753e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000110000111100110111000100;
		x2 = 32'b10000011000011100110001000101111;
		correct = 32'b00010000110000111100110111000100;
		#400; //7.723097e-29 * -4.184276e-37 = 7.723097e-29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001110110111010010100000010101;
		x2 = 32'b10000111100110100010000000001101;
		correct = 32'b01001110110111010010100000010101;
		#400; //1855195800.0 * -2.3190182e-34 = 1855195800.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001110100011111000000111010;
		x2 = 32'b01100111100101000111100100011000;
		correct = 32'b11100111100101001000011000110111;
		#400; //-4.8408496e+20 * 1.402288e+24 = -1.4027721e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000100110001011011010110100010;
		x2 = 32'b10000111100111010101010101100000;
		correct = 32'b11000100110001011011010110100010;
		#400; //-1581.676 * -2.3672913e-34 = -1581.676
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001100110011100010100000000011;
		x2 = 32'b10010110111010110110101000001100;
		correct = 32'b00010110111010110110101000011001;
		#400; //3.1763407e-31 * -3.8033223e-25 = 3.8033255e-25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110011110100000111111000001001;
		x2 = 32'b11101011011101001010101001010001;
		correct = 32'b01101011011101001010101001010001;
		#400; //9.7086804e-08 * -2.957822e+26 = 2.957822e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001110001000001100110100000;
		x2 = 32'b00010000111001001100111001001001;
		correct = 32'b11100001110001000001100110100000;
		#400; //-4.5217604e+20 * 9.0247976e-29 = -4.5217604e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100000110111100010110010111101;
		x2 = 32'b01101101000110000111110110010000;
		correct = 32'b11101101000110000111110110010000;
		#400; //1.2807503e+20 * 2.9495948e+27 = -2.9495948e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100001100110111010010110001100;
		x2 = 32'b11101101011110100001000101101000;
		correct = 32'b01101101011110100001000101101001;
		#400; //3.5889678e+20 * -4.8370185e+27 = 4.8370188e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011110101100100000001000000000;
		x2 = 32'b01111110101111001010011110100100;
		correct = 32'b11111110101111001010011110100100;
		#400; //-6.4134073e+18 * 1.2538265e+38 = -1.2538265e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011100100011100100100110110001;
		x2 = 32'b10010101010111100010101010111001;
		correct = 32'b01011100100011100100100110110001;
		#400; //3.2040377e+17 * -4.4866245e-26 = 3.2040377e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101110101010011011010110011;
		x2 = 32'b10001000101100111110011010111100;
		correct = 32'b01111101110101010011011010110011;
		#400; //3.5426197e+37 * -1.0827416e-33 = 3.5426197e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010110111000110111010001101111;
		x2 = 32'b10001000100100000011011001111011;
		correct = 32'b10010110111000110111010001101111;
		#400; //-3.6747308e-25 * -8.679493e-34 = -3.6747308e-25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110010101110010000101000010;
		x2 = 32'b11110110100000000110011111011100;
		correct = 32'b01110110100000000110011111011100;
		#400; //-3.2056855e-06 * -1.3021885e+33 = 1.3021885e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011100001011111101010101010011;
		x2 = 32'b11110101000001001011011101100000;
		correct = 32'b01110101000001001011011101100000;
		#400; //-1.979707e+17 * -1.682379e+32 = 1.682379e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100111100100001011001111001;
		x2 = 32'b01110010010010001001110100100011;
		correct = 32'b11110010010010001001110100100011;
		#400; //-0.029551731 * 3.973566e+30 = -3.973566e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011111011100101100000110000101;
		x2 = 32'b11000111110001000111010001110000;
		correct = 32'b01011111011100101100000110000101;
		#400; //1.7492409e+19 * -100584.875 = 1.7492409e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000111011111100101001010010000;
		x2 = 32'b11110101111111011010001110000110;
		correct = 32'b01110101111111011010001110000110;
		#400; //65106.562 * -6.4305066e+32 = 6.4305066e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000101001111001100100000011001;
		x2 = 32'b01010011010110001010001011101010;
		correct = 32'b11010011010110001010001011101010;
		#400; //-3020.506 * 930446200000.0 = -930446200000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001001110101010101000101010010;
		x2 = 32'b10001000110001101001000100100011;
		correct = 32'b00001010000000110111101011001101;
		#400; //5.1354358e-33 * -1.1950813e-33 = 6.330517e-33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111000101010010110010000110011;
		x2 = 32'b11101100000000110010011011011000;
		correct = 32'b11111000101010010110010000110011;
		#400; //-2.7485327e+34 * -6.342109e+26 = -2.7485327e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000001101011011001000010111101;
		x2 = 32'b01101100011001101101001100011100;
		correct = 32'b11101100011001101101001100011100;
		#400; //6.375785e-38 * 1.1161995e+27 = -1.1161995e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011001100001110110101000011010;
		x2 = 32'b11010001000111000101000100111011;
		correct = 32'b01011001100001110110101001101000;
		#400; //4764472700000000.0 * -41961107000.0 = 4764514600000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110101001100011111001010010;
		x2 = 32'b00111000111111011110011001111001;
		correct = 32'b00111110101001100010111001110100;
		#400; //0.32469422 * 0.00012106909 = 0.32457316
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001101010001101000100010011000;
		x2 = 32'b01010100110111001101100011011010;
		correct = 32'b11010100110111001101011101001101;
		#400; //208177540.0 * 7588248000000.0 = -7588039600000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011000111100101100100110000000;
		x2 = 32'b10111010111100000010011101111100;
		correct = 32'b01011000111100101100100110000000;
		#400; //2135578000000000.0 * -0.0018322314 = 2135578000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011101001001101010010001000110;
		x2 = 32'b10011011110010011001000001011001;
		correct = 32'b01011101001001101010010001000110;
		#400; //7.504875e+17 * -3.3345943e-22 = 7.504875e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111000111001011000100101111;
		x2 = 32'b00010101110101010000111100100101;
		correct = 32'b00110111000111001011000100101111;
		#400; //9.339578e-06 * 8.605391e-26 = 9.339578e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001010111000101100001010010011;
		x2 = 32'b01001001010101110111101000000101;
		correct = 32'b11001001010101110111101000000101;
		#400; //-2.1836199e-32 * 882592.3 = -882592.3
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001110101100101101011001010111;
		x2 = 32'b11110010110010010011111001111011;
		correct = 32'b01110010110010010011111001111011;
		#400; //-4.408679e-30 * -7.972099e+30 = 7.972099e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001010100110010010010110000;
		x2 = 32'b00000011001100100100001011011101;
		correct = 32'b00101001010100110010010010110000;
		#400; //4.6883233e-14 * 5.2386254e-37 = 4.6883233e-14
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101000001110111100111111001111;
		x2 = 32'b10011011110101010110010001001011;
		correct = 32'b11101000001110111100111111001111;
		#400; //-3.5476637e+24 * -3.5302707e-22 = -3.5476637e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111001010111001111101111010101;
		x2 = 32'b01011111111100010110011100000010;
		correct = 32'b11011111111100010110011100000010;
		#400; //-0.0002107465 * 3.4789749e+19 = -3.4789749e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001001001100011000110001000110;
		x2 = 32'b00001101101000010111110101101110;
		correct = 32'b10001101101000010010010010101000;
		#400; //2.1371556e-33 * 9.952587e-31 = -9.931216e-31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100110111001001001110100101110;
		x2 = 32'b01010010011101110001010101100001;
		correct = 32'b01100110111001001001110100101110;
		#400; //5.397995e+23 * 265303900000.0 = 5.397995e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001010011010011001010000111010;
		x2 = 32'b00000011001010101000001011010101;
		correct = 32'b00001010011010011001000110010000;
		#400; //1.124642e-32 * 5.0108698e-37 = 1.1245919e-32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000101011000000011001001101110;
		x2 = 32'b01101001001101001101011000010000;
		correct = 32'b11101001001101001101011000010000;
		#400; //3587.1519 * 1.3663596e+25 = -1.3663596e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110001000000000101011000111011;
		x2 = 32'b10111011101001000100010101010000;
		correct = 32'b00111011101001000100010101010100;
		#400; //1.8675468e-09 * -0.0050131455 = 0.0050131474
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001000111110001001010110010011;
		x2 = 32'b01101000000011010100111101011000;
		correct = 32'b11101000000011010100111101011000;
		#400; //-509100.6 * 2.6692692e+24 = -2.6692692e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011001111101000001110100000100;
		x2 = 32'b00110111001110010001010010110011;
		correct = 32'b10110111001110010001010010110011;
		#400; //-2.5240728e-23 * 1.1031679e-05 = -1.1031679e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111010110110001111010110100110;
		x2 = 32'b11111000110100111101011101010011;
		correct = 32'b01111000110100111101011101010011;
		#400; //-0.0016552701 * -3.4373185e+34 = 3.4373185e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101101111111000110001111011110;
		x2 = 32'b00101010101011110110000111010110;
		correct = 32'b01101101111111000110001111011110;
		#400; //9.7638693e+27 * 3.1154132e-13 = 9.7638693e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110000001011011101100101111100;
		x2 = 32'b10001111000101011011010100101101;
		correct = 32'b00110000001011011101100101111100;
		#400; //6.32461e-10 * -7.38116e-30 = 6.32461e-10
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111110101011111111000100011100;
		x2 = 32'b01011101100011111100101011001111;
		correct = 32'b01111110101011111111000100011100;
		#400; //1.1693341e+38 * 1.2951652e+18 = 1.1693341e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011110101011001010011111001;
		x2 = 32'b10111110000100110000110111001101;
		correct = 32'b00111110000100110000110111001101;
		#400; //2.3156599e-17 * -0.14360733 = 0.14360733
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001011100010010110100011101111;
		x2 = 32'b10100111010011000100111011000100;
		correct = 32'b00100111010011000100111011000100;
		#400; //-5.2928367e-32 * -2.8353386e-15 = 2.8353386e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001100101100110001011110111001;
		x2 = 32'b01011110111110110100110010001100;
		correct = 32'b11011110111110110100110010001100;
		#400; //-2.7593594e-31 * 9.054001e+18 = -9.054001e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001101010000000010101010001;
		x2 = 32'b11001000111110001010101010001101;
		correct = 32'b01001000111110001010011111101101;
		#400; //-21.002596 * -509268.4 = 509247.4
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100101110000110000000000111111;
		x2 = 32'b01001000011000000011001100011110;
		correct = 32'b01100101110000110000000000111111;
		#400; //1.1510825e+23 * 229580.47 = 1.1510825e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111011101010111010111010010101;
		x2 = 32'b10100111010000011111101110100010;
		correct = 32'b01111011101010111010111010010101;
		#400; //1.7828474e+36 * -2.692054e-15 = 1.7828474e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111100001000110111010111001110;
		x2 = 32'b01110110000111010010010000010101;
		correct = 32'b01111100001000110110101111111100;
		#400; //3.394935e+36 * 7.9679926e+32 = 3.3941383e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100100011101101101000010100110;
		x2 = 32'b11001101010010001000011011011100;
		correct = 32'b01100100011101101101000010100110;
		#400; //1.8211735e+22 * -210267580.0 = 1.8211735e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011000010110000011011111010101;
		x2 = 32'b00011111001001000011100011100100;
		correct = 32'b01011000010110000011011111010101;
		#400; //950937200000000.0 * 3.477541e-20 = 950937200000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101110100010100111101100110;
		x2 = 32'b01100000100100110111110110011101;
		correct = 32'b11100000100100110111110110011101;
		#400; //-3.6309523e-16 * 8.502259e+19 = -8.502259e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101000111110010111001110001001;
		x2 = 32'b10010010110101000110010001110110;
		correct = 32'b10101000111110010111001110001001;
		#400; //-2.7694659e-14 * -1.34038465e-27 = -2.7694659e-14
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001111101101000011001111010101;
		x2 = 32'b11010111010110110111110001100110;
		correct = 32'b01010111010110110111101011111110;
		#400; //-6046591500.0 * -241327330000000.0 = 241321300000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111010011000101111110010100001;
		x2 = 32'b01001101000010110010111111010111;
		correct = 32'b11001101000010110010111111010111;
		#400; //0.00086588605 * 145948020.0 = -145948020.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010110101100010010011110110111;
		x2 = 32'b11111010001000101100011110011011;
		correct = 32'b01111010001000101100011110011011;
		#400; //-2.8620956e-25 * -2.1130014e+35 = 2.1130014e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101111110111011011000011001100;
		x2 = 32'b00111000011101110001101110010100;
		correct = 32'b10111000011101110001110000000011;
		#400; //-4.0325288e-10 * 5.8915073e-05 = -5.8915477e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111000110100110000101110100010;
		x2 = 32'b11000001100010010110110111011011;
		correct = 32'b01000001100010010110111000010000;
		#400; //0.00010063431 * -17.17864 = 17.178741
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111101010010110011101001001;
		x2 = 32'b00011010000010011101111011010000;
		correct = 32'b10110111101010010110011101001001;
		#400; //-2.0194466e-05 * 2.8510922e-23 = -2.0194466e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000110101010101000111000101011;
		x2 = 32'b01010100001111100110010111011011;
		correct = 32'b11010100001111100110010111011011;
		#400; //21831.084 * 3271010500000.0 = -3271010500000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111111001101000010101001000101;
		x2 = 32'b11101010000100111100001001100010;
		correct = 32'b01111111001101000010101001000101;
		#400; //2.3948052e+38 * -4.465751e+25 = 2.3948052e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011101001101000011001011101111;
		x2 = 32'b11011011110100111000101011100011;
		correct = 32'b11011101000110011100000110010011;
		#400; //-8.11544e+17 * -1.19087855e+17 = -6.9245614e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110000011100110000000111001000;
		x2 = 32'b11111100110011110100010001001101;
		correct = 32'b01111100110011110100010001001101;
		#400; //-8.8405416e-10 * -8.609526e+36 = 8.609526e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100001001111011011110001010101;
		x2 = 32'b11001100111100010111010001111000;
		correct = 32'b01100001001111011011110001010101;
		#400; //2.1875034e+20 * -126591940.0 = 2.1875034e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000111001010000001000001100110;
		x2 = 32'b00100001000100000000101110011111;
		correct = 32'b10100001000100000000101110011111;
		#400; //1.2643734e-34 * 4.880448e-19 = -4.880448e-19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000000011011000000100010111;
		x2 = 32'b01111110000100001111110100100011;
		correct = 32'b11111110000100001111110100100011;
		#400; //-1.7517379e+29 * 4.81808e+37 = -4.81808e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101001101011001110110111101;
		x2 = 32'b10010001011001001000110010110110;
		correct = 32'b11111101001101011001110110111101;
		#400; //-1.5088081e+37 * -1.8029389e-28 = -1.5088081e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110010100000111000000100100110;
		x2 = 32'b10011001101110011001010110111110;
		correct = 32'b11110010100000111000000100100110;
		#400; //-5.2094294e+30 * -1.9189032e-23 = -5.2094294e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011111011011001101001100110;
		x2 = 32'b01000110000001011111100001111010;
		correct = 32'b11111011111011011001101001100110;
		#400; //-2.4674119e+36 * 8574.119 = -2.4674119e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111110011100001110101100010011;
		x2 = 32'b00111101111001110010100101011001;
		correct = 32'b01111110011100001110101100010011;
		#400; //8.0058824e+37 * 0.11287183 = 8.0058824e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010011110111000010010001001010;
		x2 = 32'b00110000101011101101111101010001;
		correct = 32'b10110000101011101101111101010001;
		#400; //-5.557159e-27 * 1.2723637e-09 = -1.2723637e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100110111111100110101100101010;
		x2 = 32'b00111011100110111101001000010001;
		correct = 32'b10111011100110111101001000010001;
		#400; //-1.7653837e-15 * 0.0047552665 = -0.0047552665
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111111000111111101000111100000;
		x2 = 32'b00100000100100000010101110011110;
		correct = 32'b01111111000111111101000111100000;
		#400; //2.1243698e+38 * 2.4423412e-19 = 2.1243698e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111000111001100001111000010;
		x2 = 32'b10010000110101110001011111010011;
		correct = 32'b00100111000111001100001111000010;
		#400; //2.175547e-15 * -8.4839254e-29 = 2.175547e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000100001010101000100001010101;
		x2 = 32'b01001001110111001001110111100011;
		correct = 32'b11001001110111001011001100110100;
		#400; //-682.1302 * 1807292.4 = -1807974.5
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111011000110000101101100111;
		x2 = 32'b10001011101110000110011001010111;
		correct = 32'b11011111011000110000101101100111;
		#400; //-1.6360283e+19 * -7.1028206e-32 = -1.6360283e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111111101001001000101110111011;
		x2 = 32'b11010101000111111100011111001101;
		correct = 32'b01010101000111111100011111001101;
		#400; //1.2855142 * -10980030000000.0 = 10980030000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010000101111111100000111010011;
		x2 = 32'b11110001100111000110001101010111;
		correct = 32'b01110001100111000110001101010111;
		#400; //-7.563485e-29 * -1.5487922e+30 = 1.5487922e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011110110111000000001110000100;
		x2 = 32'b11100001000010110101100101010010;
		correct = 32'b01100001000001000111100100110110;
		#400; //-7.92683e+18 * -1.6065835e+20 = 1.5273152e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110000100011100001101101111111;
		x2 = 32'b01001000111000111110111100101001;
		correct = 32'b11001000111000111110111100101001;
		#400; //1.0339675e-09 * 466809.28 = -466809.28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000101010000010011100000100101;
		x2 = 32'b10100101100100110100000010011011;
		correct = 32'b01000101010000010011100000100101;
		#400; //3091.509 * -2.5544213e-16 = 3091.509
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110011101110100101111011101110;
		x2 = 32'b11100000001000001001001110011010;
		correct = 32'b01110011101110100101111011101110;
		#400; //2.9531635e+31 * -4.6283045e+19 = 2.9531635e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111000100011111000100110010;
		x2 = 32'b11000000101001010111110100001011;
		correct = 32'b01000000100100110011111011100101;
		#400; //-0.5700866 * -5.171514 = 4.6014276
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100101110000010111010011111;
		x2 = 32'b00100101001010111110000100001101;
		correct = 32'b10100101001010111110000101101001;
		#400; //-1.218815e-21 * 1.4908136e-16 = -1.4908258e-16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101110111000110001101011000100;
		x2 = 32'b11101101111011101111011100001101;
		correct = 32'b01101111000011110110110001000100;
		#400; //3.5142727e+28 * -9.2445123e+27 = 4.438724e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111001011011110110000011101011;
		x2 = 32'b00001010111111000011011000100101;
		correct = 32'b10111001011011110110000011101011;
		#400; //-0.00022828921 * 2.4287084e-32 = -0.00022828921
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111010010110101001000010111;
		x2 = 32'b11001110000110010110110100111011;
		correct = 32'b11010111010010110101000111110001;
		#400; //-223553430000000.0 * -643518140.0 = -223552800000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010011100001100100100001011011;
		x2 = 32'b00001000110101101011111011000010;
		correct = 32'b01010011100001100100100001011011;
		#400; //1153479100000.0 * 1.2924503e-33 = 1153479100000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001010010111101001010010110011;
		x2 = 32'b11001011010100100001110001111010;
		correct = 32'b01001011000110100111011101001101;
		#400; //-3646764.8 * -13769850.0 = 10123085.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101010111101001101110111001111;
		x2 = 32'b00000100011110101111000010000000;
		correct = 32'b00101010111101001101110111001111;
		#400; //4.3497018e-13 * 2.9497791e-36 = 4.3497018e-13
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100101101011000011110111111;
		x2 = 32'b01000011111100011010101000001101;
		correct = 32'b11000011111100011010011100110111;
		#400; //0.022159455 * 483.32852 = -483.30637
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101010011011110000011000101;
		x2 = 32'b10100100111001101100001011000100;
		correct = 32'b00111101010011011110000011000101;
		#400; //0.050263185 * -1.00076546e-16 = 0.050263185
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100101110101011010011100001011;
		x2 = 32'b00110110100000011111100001011110;
		correct = 32'b11100101110101011010011100001011;
		#400; //-1.2611818e+23 * 3.8734133e-06 = -1.2611818e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000010110001111010010110101111;
		x2 = 32'b11111001001100111010011010111100;
		correct = 32'b01111001001100111010011010111100;
		#400; //-99.8236 * -5.830018e+34 = 5.830018e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000011001000000011110010001000;
		x2 = 32'b01001111101110010011100101100100;
		correct = 32'b11001111101110010011100101100100;
		#400; //4.708926e-37 * 6215092000.0 = -6215092000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010001001110100010001101110110;
		x2 = 32'b11010101100010001100011010101001;
		correct = 32'b01010101100010001100011010101001;
		#400; //-1.468374e-28 * -18798353000000.0 = 18798353000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011000101100010011110001101010;
		x2 = 32'b00100001110000101000011000000010;
		correct = 32'b01011000101100010011110001101010;
		#400; //1558984300000000.0 * 1.3181423e-18 = 1558984300000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010000000010011111111101001101;
		x2 = 32'b01010010110110011000010011101111;
		correct = 32'b11010010110110011000010011101111;
		#400; //-2.7215163e-29 * 467119080000.0 = -467119080000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100111010011000110010111101100;
		x2 = 32'b10001111000110000100001001011000;
		correct = 32'b01100111010011000110010111101100;
		#400; //9.652429e+23 * -7.506956e-30 = 9.652429e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111111110101010111100101111110;
		x2 = 32'b01011011001011000111101011100010;
		correct = 32'b01111111110101010111100101111110;
		#400; //nan * 4.8548807e+16 = nan
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100000000111110011111101111;
		x2 = 32'b10111001111100110001000000101110;
		correct = 32'b11110100000000111110011111101111;
		#400; //-4.1802677e+31 * -0.00046360627 = -4.1802677e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101001000110001011001111111;
		x2 = 32'b01001110011001110010011000100001;
		correct = 32'b11111101001000110001011001111111;
		#400; //-1.354881e+37 * 969508900.0 = -1.354881e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010011101100101100100001010111;
		x2 = 32'b01010111110110101101100011111000;
		correct = 32'b11010111110110111000101111000000;
		#400; //-1535730600000.0 * 481250820000000.0 = -482786540000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001100111111110010001100101110;
		x2 = 32'b01011101110100100111010011100101;
		correct = 32'b11011101110100100111010011100101;
		#400; //-3.9310144e-31 * 1.8956247e+18 = -1.8956247e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101000010110001010100100101010;
		x2 = 32'b11010010010101100101001001011011;
		correct = 32'b01010010010101100101001001011011;
		#400; //1.202709e-14 * -230126170000.0 = 230126170000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110001111000010111011100010110;
		x2 = 32'b11011011000110000111101000100001;
		correct = 32'b01011011000110000111101000100001;
		#400; //-6.5619004e-09 * -4.291848e+16 = 4.291848e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101100101010001110111010110001;
		x2 = 32'b10101100001011110100110101111101;
		correct = 32'b01101100101010001110111010110001;
		#400; //1.6338138e+27 * -2.491201e-12 = 1.6338138e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110000100010000100111101110;
		x2 = 32'b10110100101011010001010000100010;
		correct = 32'b11111110000100010000100111101110;
		#400; //-4.8197404e+37 * -3.223841e-07 = -4.8197404e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100110000000000111000100101;
		x2 = 32'b01111101101101011100111010110000;
		correct = 32'b11111101101101011100111010110000;
		#400; //-5.4585386e-12 * 3.020793e+37 = -3.020793e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111110100010001110101011101001;
		x2 = 32'b00111011100111011000011001011110;
		correct = 32'b10111110100010110110000100000010;
		#400; //-0.26741722 * 0.0048072776 = -0.2722245
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001011001110100010001100111;
		x2 = 32'b11110011100110100011111101110111;
		correct = 32'b01110011100110100011111101110111;
		#400; //-4.2477075e-38 * -2.4441557e+31 = 2.4441557e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111101010010100110101000101010;
		x2 = 32'b10001001111100000111110110010100;
		correct = 32'b10111101010010100110101000101010;
		#400; //-0.049417652 * -5.789599e-33 = -0.049417652
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110110011110011000101111010111;
		x2 = 32'b11010000100111110101000111000000;
		correct = 32'b01110110011110011000101111010111;
		#400; //1.2653498e+33 * -21383480000.0 = 1.2653498e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010001010110010111001110011100;
		x2 = 32'b00100110110101110110001110110010;
		correct = 32'b01010001010110010111001110011100;
		#400; //58371720000.0 * 1.4945644e-15 = 58371720000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001101000010110110000111011100;
		x2 = 32'b01101000010100110010010110010011;
		correct = 32'b11101000010100110010010110010011;
		#400; //4.2950476e-31 * 3.9884498e+24 = -3.9884498e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010110101001100010011101100001;
		x2 = 32'b10110000010010001110110011001110;
		correct = 32'b01010110101001100010011101100001;
		#400; //91344030000000.0 * -7.3096096e-10 = 91344030000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110110110110100101111001100;
		x2 = 32'b00010011000010010011100001010111;
		correct = 32'b00100110110110110100101111001100;
		#400; //1.5216722e-15 * 1.7319609e-27 = 1.5216722e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101110010110000111111001011101;
		x2 = 32'b01011011010101011001100100010111;
		correct = 32'b11011011010101011001100100010111;
		#400; //4.9224947e-11 * 6.0122494e+16 = -6.0122494e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010010000111001000100001111100;
		x2 = 32'b10010010110001111101010101111000;
		correct = 32'b00010011000010110000110011011011;
		#400; //4.939315e-28 * -1.261129e-27 = 1.7550605e-27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110100110110111011111111110;
		x2 = 32'b11001110010101011010011001011001;
		correct = 32'b01001110010101011010011001011001;
		#400; //-7.069899e-11 * -896112200.0 = 896112200.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101101111110001001000000100110;
		x2 = 32'b10111100110010000111001110100000;
		correct = 32'b01101101111110001001000000100110;
		#400; //9.6158184e+27 * -0.024469197 = 9.6158184e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110001011101110100010110000;
		x2 = 32'b01000001011000101100110010011011;
		correct = 32'b11111110001011101110100010110000;
		#400; //-5.8123463e+37 * 14.1749525 = -5.8123463e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101001001000111101011100110010;
		x2 = 32'b10110001001010001000001001110110;
		correct = 32'b00110001001010001000000111010010;
		#400; //-3.6379923e-14 * -2.4521376e-09 = 2.4521012e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000000110010011101111000110;
		x2 = 32'b10111011110001100010001111101010;
		correct = 32'b11110000000110010011101111000110;
		#400; //-1.8969387e+29 * -0.0060467618 = -1.8969387e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000100111001001010101010100111;
		x2 = 32'b10011011110110000011011100001001;
		correct = 32'b00011011110110000011011100001001;
		#400; //5.3759262e-36 * -3.5769768e-22 = 3.5769768e-22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001100011001011011100001010;
		x2 = 32'b10010001010110111011100110011100;
		correct = 32'b11000001100011001011011100001010;
		#400; //-17.589375 * -1.7333249e-28 = -17.589375
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011001011011001100010010010101;
		x2 = 32'b10000010010100010010110100110000;
		correct = 32'b10011001011011001100010010010101;
		#400; //-1.22406135e-23 * -1.5367863e-37 = -1.22406135e-23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001001111100110110000100010101;
		x2 = 32'b10100111001001101010100100111110;
		correct = 32'b00100111001001101010100100111110;
		#400; //5.8591418e-33 * -2.3128874e-15 = 2.3128874e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111001010010111010001110110;
		x2 = 32'b10000001100001111010100010110000;
		correct = 32'b00110111001010010111010001110110;
		#400; //1.0100301e-05 * -4.983322e-38 = 1.0100301e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001101010100011110101110110110;
		x2 = 32'b00101010110101100011111011110001;
		correct = 32'b11001101010100011110101110110110;
		#400; //-220117860.0 * 3.805771e-13 = -220117860.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000010001010101111011010111001;
		x2 = 32'b00100100100100101111111011101111;
		correct = 32'b10100100100100101111111011101111;
		#400; //1.2560433e-37 * 6.374928e-17 = -6.374928e-17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101110100110100001000101010110;
		x2 = 32'b11011000101011010100010110100001;
		correct = 32'b11101110100110100001000101010110;
		#400; //-2.3840825e+28 * -1524116500000000.0 = -2.3840825e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000101100111000110001101101;
		x2 = 32'b10111100101111100010101100111101;
		correct = 32'b01010000101100111000110001101101;
		#400; //24098597000.0 * -0.023213977 = 24098597000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111111011001011101011011101;
		x2 = 32'b10101000001110111111101101100110;
		correct = 32'b11111111111011001011101011011101;
		#400; //nan * -1.0435099e-14 = nan
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100111111101100100101101110101;
		x2 = 32'b10101111101110101100100101100101;
		correct = 32'b11100111111101100100101101110101;
		#400; //-2.3261882e+24 * -3.3976302e-10 = -2.3261882e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101111111111100001100011011101;
		x2 = 32'b01010000101111110110111100100111;
		correct = 32'b11010000101111110110111100100111;
		#400; //-4.6219997e-10 * 25693862000.0 = -25693862000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110011111110011111110101101;
		x2 = 32'b01011111111101010011100001111000;
		correct = 32'b11011111111101010011100001111000;
		#400; //4.800695e-35 * 3.534001e+19 = -3.534001e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001110110100111010001101100;
		x2 = 32'b00001100101110111110101100010011;
		correct = 32'b11100001110110100111010001101100;
		#400; //-5.037224e+20 * 2.8953392e-31 = -5.037224e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011000000110100101010101100111;
		x2 = 32'b00110110101111010111000100010011;
		correct = 32'b10110110101111010111000100010011;
		#400; //1.994715e-24 * 5.6458025e-06 = -5.6458025e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110110110011110011100101010000;
		x2 = 32'b00011000100111100111100001010101;
		correct = 32'b01110110110011110011100101010000;
		#400; //2.1014998e+33 * 4.0963547e-24 = 2.1014998e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100000010011000110001101010110;
		x2 = 32'b10101101110110000001000010101101;
		correct = 32'b01100000010011000110001101010110;
		#400; //5.891084e+19 * -2.4563762e-11 = 5.891084e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011010101011111101101100110;
		x2 = 32'b10100100010011010001111010010010;
		correct = 32'b01101011010101011111101101100110;
		#400; //2.586884e+26 * -4.4478183e-17 = 2.586884e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000011001111001010001000111011;
		x2 = 32'b10010101110001011000101000101111;
		correct = 32'b00010101110001011000101000101111;
		#400; //5.5434466e-37 * -7.978568e-26 = 7.978568e-26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111000001101100111000001101101;
		x2 = 32'b00101101100101100101001111010000;
		correct = 32'b10111000001101100111000001110010;
		#400; //-4.3496886e-05 * 1.7090246e-11 = -4.3496904e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011000011111000000111101010011;
		x2 = 32'b00000111111010011011100010110100;
		correct = 32'b11011000011111000000111101010011;
		#400; //-1108571000000000.0 * 3.5166502e-34 = -1108571000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000101110000001000011100011010;
		x2 = 32'b10001010000001100001010001001000;
		correct = 32'b00001010000001011011010000000100;
		#400; //-1.8105222e-35 * -6.45568e-33 = 6.437574e-33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010010110011000001110111111010;
		x2 = 32'b01001111110100011001011001111110;
		correct = 32'b01010010110010001101011110100000;
		#400; //438338130000.0 * 7032601600.0 = 431305520000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100101100000010100100001101;
		x2 = 32'b00110100011000111001110100011110;
		correct = 32'b11111100101100000010100100001101;
		#400; //-7.317415e+36 * 2.1198181e-07 = -7.317415e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011100111011010011001000100010;
		x2 = 32'b01011110111001001111010100000111;
		correct = 32'b11011110110101100010000111100101;
		#400; //5.3411753e+17 * 8.24905e+18 = -7.714933e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001000101011010110101001101101;
		x2 = 32'b00001110011011110101011110111110;
		correct = 32'b10001110011011110100001000010001;
		#400; //1.0437079e-33 * 2.950127e-30 = -2.9490834e-30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110011000011100101111101010110;
		x2 = 32'b11100001111101111111111010001101;
		correct = 32'b11110011000011100101111101010110;
		#400; //-1.1279904e+31 * -5.71836e+20 = -1.1279904e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100110100110011010001000111011;
		x2 = 32'b11001111001110111110110111011000;
		correct = 32'b01100110100110011010001000111011;
		#400; //3.6275735e+23 * -3152926700.0 = 3.6275735e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001101101001001101000110101;
		x2 = 32'b10001100011010000100111110101010;
		correct = 32'b01111001101101001001101000110101;
		#400; //1.1721764e+35 * -1.7896603e-31 = 1.1721764e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111000100011000000011101011010;
		x2 = 32'b01100010110000110001110101110011;
		correct = 32'b01111000100011000000011101011010;
		#400; //2.2720958e+34 * 1.7996186e+21 = 2.2720958e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001111111100000001011000011100;
		x2 = 32'b11000011010100001110100101000000;
		correct = 32'b11001111111100000001011000011100;
		#400; //-8055961600.0 * -208.91113 = -8055961600.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100110000010011110011110010;
		x2 = 32'b01111000111001101100001111011001;
		correct = 32'b11111000111001111000010100010110;
		#400; //-1.2247918e+32 * 3.7443767e+34 = -3.7566246e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111011100010110011010101011011;
		x2 = 32'b10100010010111001001110000001101;
		correct = 32'b00111011100010110011010101011011;
		#400; //0.004248304 * -2.9898172e-18 = 0.004248304
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110010100011100101001111110;
		x2 = 32'b10011010100110110111110011000111;
		correct = 32'b11111110010100011100101001111110;
		#400; //-6.9715013e+37 * -6.4308086e-23 = -6.9715013e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110011001100101000111001000000;
		x2 = 32'b00001100101011001010110000011101;
		correct = 32'b00110011001100101000111001000000;
		#400; //4.157323e-08 * 2.6604383e-31 = 4.157323e-08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010111100010011010000001110110;
		x2 = 32'b10000000000000000110100001111111;
		correct = 32'b01010111100010011010000001110110;
		#400; //302644530000000.0 * -3.7486e-41 = 302644530000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001111000111011000010110110110;
		x2 = 32'b10100000101011100000111000001000;
		correct = 32'b00100000101011100000111000001000;
		#400; //-7.7664494e-30 * -2.9486032e-19 = 2.9486032e-19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000100110010101111001010111000;
		x2 = 32'b01100111000100010101100111001110;
		correct = 32'b11100111000100010101100111001110;
		#400; //4.7712874e-36 * 6.8639974e+23 = -6.8639974e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001000101111110001010111011110;
		x2 = 32'b01110101101011010111101100011100;
		correct = 32'b11110101101011010111101100011100;
		#400; //391342.94 * 4.3982632e+32 = -4.3982632e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111000010110001001110000011000;
		x2 = 32'b00110110001011010001110010111000;
		correct = 32'b10111000011000110110110111100100;
		#400; //-5.1643787e-05 * 2.5795725e-06 = -5.422336e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110110101111000111001111100;
		x2 = 32'b11001001111000100011111100011001;
		correct = 32'b01001001111000100011111100011001;
		#400; //1.4957242e-15 * -1853411.1 = 1853411.1
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011100010010001101100100100010;
		x2 = 32'b01110011100011001000001111011100;
		correct = 32'b11110011100011001000001111011100;
		#400; //2.2613494e+17 * 2.2265503e+31 = -2.2265503e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010101011111000001000000100101;
		x2 = 32'b11111010101111000010010000100010;
		correct = 32'b01111010101111000010010000100010;
		#400; //17321642000000.0 * -4.8844233e+35 = 4.8844233e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011100001111011101011010110;
		x2 = 32'b11101111101110001000001001111110;
		correct = 32'b11111011100001111011101011010101;
		#400; //-1.4094991e+36 * -1.1420599e+29 = -1.409499e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011111001001001000111111111110;
		x2 = 32'b11100111101001101101000111000011;
		correct = 32'b01100111101001101101001000010101;
		#400; //1.1857976e+19 * -1.5755645e+24 = 1.5755763e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110100000111101010111101111;
		x2 = 32'b11111001110010110110010010110000;
		correct = 32'b01111001110010110110010010110000;
		#400; //-3.9290094e-06 * -1.3200981e+35 = 1.3200981e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100010110101010000110001111;
		x2 = 32'b10011011111000001100100110010100;
		correct = 32'b10101100010110101010000110001111;
		#400; //-3.1069346e-12 * -3.7187958e-22 = -3.1069346e-12
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001110000001000011110001001;
		x2 = 32'b01000110110101111010100001101011;
		correct = 32'b11000110110101111010100001101011;
		#400; //-7.0724144e-38 * 27604.209 = -27604.209
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111000110011001110110110011111;
		x2 = 32'b00001010101110101001001110101010;
		correct = 32'b10111000110011001110110110011111;
		#400; //-9.7717384e-05 * 1.7966694e-32 = -9.7717384e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011101000101001110110010111110;
		x2 = 32'b10011110101110100100111001001010;
		correct = 32'b01011101000101001110110010111110;
		#400; //6.7069756e+17 * -1.9725896e-20 = 6.7069756e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001101100100101000000001110011;
		x2 = 32'b11010111000111100011010100011011;
		correct = 32'b01010111000111100011010100011011;
		#400; //-9.028868e-31 * -173950920000000.0 = 173950920000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011010101111001010001110100000;
		x2 = 32'b00011011111100001010100100100010;
		correct = 32'b01011010101111001010001110100000;
		#400; //2.6548602e+16 * 3.981397e-22 = 2.6548602e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110100100110000100101110000;
		x2 = 32'b10111010011011100000011100101001;
		correct = 32'b00111010011011100000011100101001;
		#400; //1.0202732e-15 * -0.00090800464 = 0.00090800464
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101111101000000000001000010110;
		x2 = 32'b01011000101110000100010000010111;
		correct = 32'b11101111101000000000001000010110;
		#400; //-9.904025e+28 * 1620820700000000.0 = -9.904025e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111000101101000100001101001;
		x2 = 32'b11110111110010001111011110100100;
		correct = 32'b01110111110010001111011110100100;
		#400; //-8.972457e-06 * -8.152204e+33 = 8.152204e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100000110110100011111001110111;
		x2 = 32'b10011010011000111011011110010110;
		correct = 32'b11100000110110100011111001110111;
		#400; //-1.258091e+20 * -4.70908e-23 = -1.258091e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100101011001000101100001010110;
		x2 = 32'b10100111000001000000000000101110;
		correct = 32'b01100101011001000101100001010110;
		#400; //6.7395567e+22 * -1.8318777e-15 = 6.7395567e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100110011000101001111011001000;
		x2 = 32'b10111100010110110100001000001000;
		correct = 32'b01100110011000101001111011001000;
		#400; //2.6754596e+23 * -0.013382442 = 2.6754596e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110011110100101010111010011110;
		x2 = 32'b10010010111111001010100000011101;
		correct = 32'b11110011110100101010111010011110;
		#400; //-3.338391e+31 * -1.5944879e-27 = -3.338391e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011101001010100101100001111;
		x2 = 32'b00101111000011001000010011000011;
		correct = 32'b01101011101001010100101100001111;
		#400; //3.9965443e+26 * 1.2780092e-10 = 3.9965443e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111010000101111011101101101;
		x2 = 32'b01010011100110111001101100011000;
		correct = 32'b11011111010000101111011101101110;
		#400; //-1.4048817e+19 * 1336644000000.0 = -1.4048819e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000011101001101000111101100;
		x2 = 32'b00011111011000111100000101010010;
		correct = 32'b10011111011000111100000101010010;
		#400; //4.8282233e-29 * 4.822903e-20 = -4.822903e-20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101100000101110010000010100011;
		x2 = 32'b11111100100001011111010010100100;
		correct = 32'b01111100100001011111010010100100;
		#400; //2.1476508e-12 * -5.564299e+36 = 5.564299e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100011101010100101001001100101;
		x2 = 32'b01001001100001110000010001011111;
		correct = 32'b11001001100001110000010001011111;
		#400; //-1.8466332e-17 * 1106059.9 = -1106059.9
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111111001100101111100100110;
		x2 = 32'b10100010011100110111000010000100;
		correct = 32'b10111111111001100101111100100110;
		#400; //-1.7997787 * -3.2992206e-18 = -1.7997787
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101100010010101101001000010111;
		x2 = 32'b11011100110111001000100100110110;
		correct = 32'b01011100110111001000100100110110;
		#400; //2.882255e-12 * -4.9660288e+17 = 4.9660288e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100110001100111100111100100101;
		x2 = 32'b11101010100111011001011100001011;
		correct = 32'b01101010100111010011110100100011;
		#400; //-2.1228119e+23 * -9.525732e+25 = 9.504503e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111010000101011110010011010100;
		x2 = 32'b11000110100011000110110111010000;
		correct = 32'b01000110100011000110110111010000;
		#400; //-0.0005717997 * -17974.906 = 17974.906
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110000110101111001100011000010;
		x2 = 32'b01110101010100011000000001011100;
		correct = 32'b11110101010100011000000001011100;
		#400; //1.5686725e-09 * 2.6557458e+32 = -2.6557458e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110001000111110000010000101110;
		x2 = 32'b11000100100100111001111010000110;
		correct = 32'b01110001000111110000010000101110;
		#400; //7.874107e+29 * -1180.9539 = 7.874107e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010100001011011110010101110;
		x2 = 32'b00110110000011011100010011001110;
		correct = 32'b10110110000011011100010011001111;
		#400; //-2.375647e-13 * 2.1125193e-06 = -2.1125195e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010010011100101101101111111010;
		x2 = 32'b11000001010001010011111111001011;
		correct = 32'b11010010011100101101101111111010;
		#400; //-260768170000.0 * -12.328074 = -260768170000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000000110010010110101010000010;
		x2 = 32'b10110101100001111000100001110010;
		correct = 32'b01000000110010010110101010000100;
		#400; //6.2942514 * -1.0097995e-06 = 6.2942524
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000111110101011001010100001010;
		x2 = 32'b10101110101001101110011010101000;
		correct = 32'b01000111110101011001010100001010;
		#400; //109354.08 * -7.589779e-11 = 109354.08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001101001010011101011000001101;
		x2 = 32'b10001011011101100111011101010100;
		correct = 32'b01001101001010011101011000001101;
		#400; //178086100.0 * -4.746765e-32 = 178086100.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001100110110010000111100100010;
		x2 = 32'b11110100110110010101011101101110;
		correct = 32'b01110100110110010101011101101110;
		#400; //3.3443252e-31 * -1.3775656e+32 = 1.3775656e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101011101100101111001011111101;
		x2 = 32'b11111100111101010001100001000101;
		correct = 32'b01111100111101010001100001000101;
		#400; //1.2715103e-12 * -1.018084e+37 = 1.018084e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100010101111110011110101101100;
		x2 = 32'b11000011110100010100111011100111;
		correct = 32'b01100010101111110011110101101100;
		#400; //1.763877e+21 * -418.61642 = 1.763877e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000100111010000100101000111100;
		x2 = 32'b01011111001110000011000110101001;
		correct = 32'b11011111001110000011000110101001;
		#400; //-5.461111e-36 * 1.3272575e+19 = -1.3272575e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101111110100101110011111111001;
		x2 = 32'b00111010010111011001111011000110;
		correct = 32'b01101111110100101110011111111001;
		#400; //1.3054458e+29 * 0.000845414 = 1.3054458e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011101100110001011011101110011;
		x2 = 32'b10001001010010011110010101110110;
		correct = 32'b00011101100110001011011101110011;
		#400; //4.0423747e-21 * -2.4302387e-33 = 4.0423747e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011001100000010111101010010111;
		x2 = 32'b00001100100000001100101011111101;
		correct = 32'b00011001100000010111101010010111;
		#400; //1.3387801e-23 * 1.9843692e-31 = 1.3387801e-23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101000000110100010100101101;
		x2 = 32'b00100010011100101010101111000011;
		correct = 32'b10100010011100101010101111000011;
		#400; //6.172296e-36 * 3.2888046e-18 = -3.2888046e-18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001111010100111010100000100;
		x2 = 32'b10000010010101101111111110101001;
		correct = 32'b11100001111010100111010100000100;
		#400; //-5.4062125e+20 * -1.5795608e-37 = -5.4062125e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011101001011011101100010011111;
		x2 = 32'b11000100110001011011101111011010;
		correct = 32'b01000100110001011011101111011010;
		#400; //-2.300835e-21 * -1581.8704 = 1581.8704
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100111011101010100111100110100;
		x2 = 32'b11010101011111111111001110010100;
		correct = 32'b11100111011101010100111100110100;
		#400; //-1.1584408e+24 * -17588852000000.0 = -1.1584408e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010000000000111101111101101110;
		x2 = 32'b00110011000110010110110000101110;
		correct = 32'b10110011000110010110110000101110;
		#400; //-2.600732e-29 * 3.5721477e-08 = -3.5721477e-08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010011101001011110101000110000;
		x2 = 32'b00011010110000101111110110110001;
		correct = 32'b01010011101001011110101000110000;
		#400; //1425197200000.0 * 8.064638e-23 = 1425197200000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000111000000001111011010001010;
		x2 = 32'b00110111101111111100100011000001;
		correct = 32'b10110111101111111100100011000001;
		#400; //9.702101e-35 * 2.2862458e-05 = -2.2862458e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011011010001100100101011101100;
		x2 = 32'b10100011111011010111111001011110;
		correct = 32'b01011011010001100100101011101100;
		#400; //5.5814423e+16 * -2.574911e-17 = 5.5814423e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001000100001010101010000000111;
		x2 = 32'b10000001110000001100110100010010;
		correct = 32'b11001000100001010101010000000111;
		#400; //-273056.22 * -7.082392e-38 = -273056.22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011011000001100010110011111001;
		x2 = 32'b11100001100100000001111000111110;
		correct = 32'b01100001100100000010001001101111;
		#400; //3.7767095e+16 * -3.323138e+20 = 3.3235154e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100101111001010110000101110111;
		x2 = 32'b10110010101010110101101111010001;
		correct = 32'b11100101111001010110000101110111;
		#400; //-1.3540248e+23 * -1.9948773e-08 = -1.3540248e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000111101101111010101000110010;
		x2 = 32'b11001110000110111010110100011001;
		correct = 32'b01001110000110111010110100011001;
		#400; //-2.7634811e-34 * -652953150.0 = 652953150.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101101101111010000011110001001;
		x2 = 32'b10010011001001000000010001110111;
		correct = 32'b00101101101111010000011110001001;
		#400; //2.1490159e-11 * -2.0701911e-27 = 2.1490159e-11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101101011000111011011000011;
		x2 = 32'b00001110001111111010101011100001;
		correct = 32'b01111101101011000111011011000011;
		#400; //2.8655483e+37 * 2.3624843e-30 = 2.8655483e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011010010110000111101110000;
		x2 = 32'b11010111100111111110011001110100;
		correct = 32'b01010111100111111110011001110100;
		#400; //1.1007921e-17 * -351624270000000.0 = 351624270000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010011000111000001000110101;
		x2 = 32'b01010011110110101100001110101001;
		correct = 32'b11010011110110101100001110101001;
		#400; //-2.0206825e-13 * 1879171000000.0 = -1879171000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011011000101101011011010011000;
		x2 = 32'b00011011101111000010001011000011;
		correct = 32'b10011011011000011000111011101110;
		#400; //1.2466708e-22 * 3.1124455e-22 = -1.8657747e-22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100100110000101110111011100;
		x2 = 32'b00100101111001001101111101101111;
		correct = 32'b00111100100110000101110111011100;
		#400; //0.018599443 * 3.97031e-16 = 0.018599443
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001110000111100101101010001000;
		x2 = 32'b11100001001111111101001011000000;
		correct = 32'b01100001001111111101001011000000;
		#400; //-664183300.0 * -2.2115714e+20 = 2.2115714e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011110001010100001011010010110;
		x2 = 32'b11110001001110010000100100101100;
		correct = 32'b01110001001110010000100100101100;
		#400; //-3.064037e+18 * -9.1625304e+29 = 9.1625304e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110010110010101110101110001100;
		x2 = 32'b01111111000100011011100110100000;
		correct = 32'b11111111000100011011100110100000;
		#400; //-8.0384935e+30 * 1.9370188e+38 = -1.9370188e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100011100100101000001001111000;
		x2 = 32'b11011000011010100101011000111000;
		correct = 32'b01011000011010100101011000111000;
		#400; //-1.5884607e-17 * -1030624100000000.0 = 1030624100000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111010001001110011110100000;
		x2 = 32'b00101111100101001100100011011110;
		correct = 32'b11011111010001001110011110100000;
		#400; //-1.4188485e+19 * 2.7063768e-10 = -1.4188485e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001110110000001101001011011;
		x2 = 32'b11000101100110101111101110100011;
		correct = 32'b01000101100110101111101110100011;
		#400; //9.596899e-14 * -4959.4546 = 4959.4546
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101110101001011000111010001101;
		x2 = 32'b01110000010110110011011101101000;
		correct = 32'b11110000010001101000010110010110;
		#400; //2.561868e+28 * 2.713768e+29 = -2.4575811e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111001111011000101100101010;
		x2 = 32'b01011001110101001111110111101110;
		correct = 32'b11011001110101001111110111101110;
		#400; //-1.12976795e-05 * 7493986700000000.0 = -7493986700000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001001110011000101110011010111;
		x2 = 32'b01011001111001001111110011010000;
		correct = 32'b11011001111001001111110011010000;
		#400; //-4.919852e-33 * 8056783000000000.0 = -8056783000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010000111111001110111101100011;
		x2 = 32'b11000110000001100011011100101111;
		correct = 32'b11010000111111001110111101011111;
		#400; //-33948375000.0 * -8589.796 = -33948367000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110100010100011000111101011001;
		x2 = 32'b10010000010100100101010011010111;
		correct = 32'b10110100010100011000111101011001;
		#400; //-1.9516791e-07 * -4.1480556e-29 = -1.9516791e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111001100101001010100110001011;
		x2 = 32'b00100000101110010011011010010011;
		correct = 32'b10111001100101001010100110001011;
		#400; //-0.0002835508 * 3.1376333e-19 = -0.0002835508
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011111111000010000111011101110;
		x2 = 32'b00011001011001000000111111100001;
		correct = 32'b01011111111000010000111011101110;
		#400; //3.2434322e+19 * 1.17905304e-23 = 3.2434322e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100100010001011100011011011;
		x2 = 32'b10111101000000010000011010110000;
		correct = 32'b00111101000000010000011010110000;
		#400; //-1.3805403e-26 * -0.03150052 = 0.03150052
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100100001001011000000010011111;
		x2 = 32'b01110100011101011101010111111100;
		correct = 32'b11110100011101011101010111111100;
		#400; //-3.5887618e-17 * 7.79085e+31 = -7.79085e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001100100111110010111000100010;
		x2 = 32'b01011010110011101111111001101011;
		correct = 32'b11011010110011101111111001101011;
		#400; //-2.4525594e-31 * 2.913179e+16 = -2.913179e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100100011001010111000000011100;
		x2 = 32'b01110011010011011010110101010001;
		correct = 32'b11110011010011011010110101010001;
		#400; //4.975142e-17 * 1.6295412e+31 = -1.6295412e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100101111110100000110000001100;
		x2 = 32'b10111101101000011100100100000110;
		correct = 32'b11100101111110100000110000001100;
		#400; //-1.4760173e+23 * -0.0789967 = -1.4760173e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110100011111100101101111011;
		x2 = 32'b01001001101111100100101011110011;
		correct = 32'b11111110100011111100101101111011;
		#400; //-9.556807e+37 * 1558878.4 = -9.556807e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011000101110000001000010111100;
		x2 = 32'b11111111010101110010010001111111;
		correct = 32'b01111111010101110010010001111111;
		#400; //4.7579783e-24 * -2.8597352e+38 = 2.8597352e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101011000101101101011011010;
		x2 = 32'b11100101110100111001001010001000;
		correct = 32'b01100101110100111001001010001000;
		#400; //0.055384494 * -1.2489029e+23 = 1.2489029e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101001101111100001110011000000;
		x2 = 32'b11100001111011011101111100011011;
		correct = 32'b01100001111011011101111100011011;
		#400; //-8.442682e-14 * -5.4849435e+20 = 5.4849435e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001000100101111110110110100;
		x2 = 32'b00011010101101111100011001110111;
		correct = 32'b01111001000100101111110110110100;
		#400; //4.7701316e+34 * 7.6007663e-23 = 4.7701316e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010100100101000101001000100011;
		x2 = 32'b10100000111000000110100100001000;
		correct = 32'b00100000111000000110100100001001;
		#400; //1.4976578e-26 * -3.801658e-19 = 3.8016582e-19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100011110100011001010101000101;
		x2 = 32'b11001001000001100101101000101110;
		correct = 32'b01001001000001100101101000101110;
		#400; //-2.2723044e-17 * -550306.9 = 550306.9
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011001010111001100100101011101;
		x2 = 32'b11011110011110101110110100010010;
		correct = 32'b01011110011110101110110100010010;
		#400; //-1.14143984e-23 * -4.520282e+18 = 4.520282e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001000011010110110011001111001;
		x2 = 32'b01011101100110111100010111010001;
		correct = 32'b11011101100110111100010111010001;
		#400; //-7.0838196e-34 * 1.4030759e+18 = -1.4030759e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000000101010100111100111001100;
		x2 = 32'b00111011010100011010110011011101;
		correct = 32'b10111011010100011010110011011101;
		#400; //1.5655727e-38 * 0.0031993904 = -0.0031993904
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111110011110000000110100110001;
		x2 = 32'b00111010011001100001000010110101;
		correct = 32'b01111110011110000000110100110001;
		#400; //8.242926e+37 * 0.0008776293 = 8.242926e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100100011001010010101000111010;
		x2 = 32'b00001100011000100110110011010010;
		correct = 32'b11100100011001010010101000111010;
		#400; //-1.6909389e+22 * 1.7443154e-31 = -1.6909389e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100100110111001111001101010;
		x2 = 32'b10001100110010001001110010011110;
		correct = 32'b00111100100110111001111001101010;
		#400; //0.018996436 * -3.090914e-31 = 0.018996436
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110001010100010011100111000001;
		x2 = 32'b11101001010110011011011011010101;
		correct = 32'b01101001010110011011011011010101;
		#400; //-3.0446332e-09 * -1.6450019e+25 = 1.6450019e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000000001111000010011100011001;
		x2 = 32'b01010000000000101001000100000011;
		correct = 32'b11010000000000101001000100000011;
		#400; //-5.524155e-39 * 8762166000.0 = -8762166000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110111010010001010100011001100;
		x2 = 32'b01010011100101111101000001010011;
		correct = 32'b11110111010010001010100011001100;
		#400; //-4.0698554e+33 * 1304070300000.0 = -4.0698554e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011100101101101110100111100;
		x2 = 32'b10110101001110011110011111001110;
		correct = 32'b01001011100101101101110100111100;
		#400; //19774072.0 * -6.925519e-07 = 19774072.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001110010110001101100100010110;
		x2 = 32'b11011101011111111001100000001001;
		correct = 32'b01011101011111111001100000001001;
		#400; //-2.6728579e-30 * -1.15109254e+18 = 1.15109254e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001101000001000000000111111010;
		x2 = 32'b00010011001101001101101110001100;
		correct = 32'b10010011001101001101001101001100;
		#400; //4.067802e-31 * 2.2827439e-27 = -2.2823371e-27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111101000011000111100011111;
		x2 = 32'b00001100110000101001100101011100;
		correct = 32'b00110111101000011000111100011111;
		#400; //1.9259342e-05 * 2.9982733e-31 = 1.9259342e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110110001001101000111100011110;
		x2 = 32'b11011001110001000000111000100001;
		correct = 32'b01110110001001101000111100011110;
		#400; //8.445547e+32 * -6898079000000000.0 = 8.445547e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001001111010110100101100010001;
		x2 = 32'b11001110000001101100011010010010;
		correct = 32'b01001110000001110011110000111000;
		#400; //1927522.1 * -565290100.0 = 567217660.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111011000000101010100110110100;
		x2 = 32'b11001111010010010101000001000110;
		correct = 32'b01001111010010010101000001000110;
		#400; //-0.0019937577 * -3377481200.0 = 3377481200.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101110011011000101000000111110;
		x2 = 32'b01111000011001000000001111100010;
		correct = 32'b11111000011001000000001111100010;
		#400; //5.3731457e-11 * 1.8498788e+34 = -1.8498788e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000101110100110000110000001101;
		x2 = 32'b00111111111011000101010010111111;
		correct = 32'b01000101110100101111110101001000;
		#400; //6753.5063 * 1.8463362 = 6751.66
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011100000111011101111001001111;
		x2 = 32'b11110000011011101111101100110001;
		correct = 32'b01110000011011101111101100110001;
		#400; //5.223427e-22 * -2.9584442e+29 = 2.9584442e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100011111011101011001000000;
		x2 = 32'b00110101011101010000010011010100;
		correct = 32'b11010100011111011101011001000000;
		#400; //-4360885000000.0 * 9.127664e-07 = -4360885000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110010010100011011111011010111;
		x2 = 32'b11011010000010000110001010001101;
		correct = 32'b11110010010100011011111011010111;
		#400; //-4.154437e+30 * -9597239000000000.0 = -4.154437e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011011001010010000001110101111;
		x2 = 32'b00000000100000111100010101111010;
		correct = 32'b01011011001010010000001110101111;
		#400; //4.757332e+16 * 1.2101291e-38 = 4.757332e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000010010100111111001010011;
		x2 = 32'b10000111110011010100011111001101;
		correct = 32'b10011000010010100111111001010011;
		#400; //-2.6171666e-24 * -3.0887172e-34 = -2.6171666e-24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001000010110100010101111000011;
		x2 = 32'b01110111010100100111010100100101;
		correct = 32'b11110111010100100111010100100101;
		#400; //-223407.05 * 4.2685872e+33 = -4.2685872e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100110110001101110100001111011;
		x2 = 32'b01010100110000011010100101111101;
		correct = 32'b11100110110001101110100001111011;
		#400; //-4.6965854e+23 * 6654178000000.0 = -4.6965854e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101001111101111000011110101;
		x2 = 32'b01010100100111011100101111110001;
		correct = 32'b11010100100111011100101111110001;
		#400; //-1.6561512e-16 * 5421851500000.0 = -5421851500000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110011011111011100001110101010;
		x2 = 32'b10000000011100101001111011011101;
		correct = 32'b01110011011111011100001110101010;
		#400; //2.010528e+31 * -1.0526236e-38 = 2.010528e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111011110000110011101001011110;
		x2 = 32'b11111100110110101001101101010100;
		correct = 32'b01111101000001011011010011110110;
		#400; //2.0273634e+36 * -9.080569e+36 = 1.1107933e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000000000110110001011000010111;
		x2 = 32'b11001010011111000001100011010001;
		correct = 32'b01001010011111000001100011010001;
		#400; //2.487483e-39 * -4130356.2 = 4130356.2
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010111001111101100001000000011;
		x2 = 32'b01100100101001000110110101001011;
		correct = 32'b11100100101001000110110101001011;
		#400; //-6.163719e-25 * 2.4265131e+22 = -2.4265131e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011110011101100000001111111101;
		x2 = 32'b00000011000110110010111101000110;
		correct = 32'b10011110011101100000001111111101;
		#400; //-1.3023956e-20 * 4.5604673e-37 = -1.3023956e-20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001001011110101000110110001010;
		x2 = 32'b11101000101010111011100001000000;
		correct = 32'b01101000101010111011100001000000;
		#400; //-1026264.6 * -6.487388e+24 = 6.487388e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111001010010000100001110111;
		x2 = 32'b00001001101011001011111001111100;
		correct = 32'b11011111001010010000100001110111;
		#400; //-1.2180116e+19 * 4.1586624e-33 = -1.2180116e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100101110000101001101100100;
		x2 = 32'b00100100101101011001100100001111;
		correct = 32'b00111100101110000101001101100100;
		#400; //0.022500701 * 7.875553e-17 = 0.022500701
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111000101000111011001111011100;
		x2 = 32'b10100101101110000010101111111001;
		correct = 32'b11111000101000111011001111011100;
		#400; //-2.6562262e+34 * -3.194871e-16 = -2.6562262e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011100100000110100011000110110;
		x2 = 32'b00110110110110011100011001101001;
		correct = 32'b10110110110110011100011001101001;
		#400; //8.687002e-22 * 6.490202e-06 = -6.490202e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111000001000110011000001010;
		x2 = 32'b10110001101110001110101101000110;
		correct = 32'b00110111000001000111110100100111;
		#400; //7.891571e-06 * -5.3818523e-09 = 7.896952e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010001111001101000010100010010;
		x2 = 32'b10100010110011010101010101011110;
		correct = 32'b11010001111001101000010100010010;
		#400; //-123759380000.0 * -5.5655747e-18 = -123759380000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110100111010110000110011000;
		x2 = 32'b00111110011111101100100100101010;
		correct = 32'b11111110100111010110000110011000;
		#400; //-1.0459777e+38 * 0.24881425 = -1.0459777e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110010111001011111101000101;
		x2 = 32'b11001010010010000000001001000111;
		correct = 32'b01001010010010000000001001000111;
		#400; //-3.2893888e-06 * -3276945.8 = 3276945.8
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101100001010011100011101100;
		x2 = 32'b10111100100110111111000101100001;
		correct = 32'b11111101100001010011100011101100;
		#400; //-2.213536e+37 * -0.019035997 = -2.213536e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001000001101100111111001110100;
		x2 = 32'b10110001110010111011101100001111;
		correct = 32'b01001000001101100111111001110100;
		#400; //186873.81 * -5.9293437e-09 = 186873.81
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001111101101100001100110110010;
		x2 = 32'b01111010011110010110100110000000;
		correct = 32'b11111010011110010110100110000000;
		#400; //-1.7956483e-29 * 3.2375543e+35 = -3.2375543e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110100110111111000101011011;
		x2 = 32'b10110011101101110001000111110010;
		correct = 32'b00111110100110111111000101011110;
		#400; //0.30457577 * -8.524866e-08 = 0.30457586
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111001111010111010101001001010;
		x2 = 32'b01001000011100100000000110000111;
		correct = 32'b11001000011100100000000110000111;
		#400; //-0.00044949568 * 247814.11 = -247814.11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100000100110100001010010001;
		x2 = 32'b01011011001000100001011010000001;
		correct = 32'b11011011001000100001011010000001;
		#400; //-2.0926908e-12 * 4.562369e+16 = -4.562369e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110010000100001010111001101010;
		x2 = 32'b01110100111100111001111010111011;
		correct = 32'b11110100111100111001111010111011;
		#400; //-8.42156e-09 * 1.5441255e+32 = -1.5441255e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101111100001011011111110100110;
		x2 = 32'b01000110100001011110111101011001;
		correct = 32'b11101111100001011011111110100110;
		#400; //-8.278639e+28 * 17143.674 = -8.278639e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111001011001010000100000110;
		x2 = 32'b10001101111010010001110110001110;
		correct = 32'b10111111001011001010000100000110;
		#400; //-0.674332 * -1.4366849e-30 = -0.674332
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001011011001011011010011100111;
		x2 = 32'b10000101010011110010111001110011;
		correct = 32'b11001011011001011011010011100111;
		#400; //-15054055.0 * -9.7416246e-36 = -15054055.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111000100100000100101110111100;
		x2 = 32'b11100011010011111110010001000010;
		correct = 32'b01100011010011111110010001000010;
		#400; //-6.880562e-05 * -3.8349237e+21 = 3.8349237e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110001101011011000011011100;
		x2 = 32'b00100100001011011111110001001001;
		correct = 32'b10110110001101011011000011011100;
		#400; //-2.7074047e-06 * 3.772709e-17 = -2.7074047e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100010110011000011000101001000;
		x2 = 32'b10011110011011111110011100010010;
		correct = 32'b01100010110011000011000101001000;
		#400; //1.8833434e+21 * -1.2700339e-20 = 1.8833434e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010010101110111101011010101111;
		x2 = 32'b00110011011010001000011110011101;
		correct = 32'b10110011011010001000011110011101;
		#400; //-1.1854283e-27 * 5.414005e-08 = -5.414005e-08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101001100111110000000101011;
		x2 = 32'b11011001100101000100110001100010;
		correct = 32'b01110101001100111110000000101011;
		#400; //2.2801948e+32 * -5217785000000000.0 = 2.2801948e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010010101110101111000000101011;
		x2 = 32'b01110111111010010011000010010011;
		correct = 32'b11110111111010010011000010010011;
		#400; //1.1797456e-27 * 9.4593e+33 = -9.4593e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011111111010101110100100000;
		x2 = 32'b01010110010100000011110011110111;
		correct = 32'b11010110010100000011110011110111;
		#400; //-1.4891384e-36 * 57240065000000.0 = -57240065000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110011001011000010001010001110;
		x2 = 32'b10000010110110110110001000101110;
		correct = 32'b10110011001011000010001010001110;
		#400; //-4.0078298e-08 * -3.223551e-37 = -4.0078298e-08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000001111110111110111101000011;
		x2 = 32'b01100001111101001100001011000001;
		correct = 32'b11100001111101001100001011000001;
		#400; //9.254616e-38 * 5.6437988e+20 = -5.6437988e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101101111000000010100011101;
		x2 = 32'b10100001111110011110011100000000;
		correct = 32'b00100001111110011110011100000000;
		#400; //1.7681313e-35 * -1.6934042e-18 = 1.6934042e-18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011011000000110100101110111;
		x2 = 32'b11111100010110101011000000000001;
		correct = 32'b01111100001000101001010110100011;
		#400; //-1.1652136e+36 * -4.541962e+36 = 3.3767483e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000010011100001010100010110001;
		x2 = 32'b01011000011001001000000100100110;
		correct = 32'b11011000011001001000000100100110;
		#400; //-1.7680827e-37 * 1004973360000000.0 = -1004973360000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100100000100010110111110000110;
		x2 = 32'b11110101110000001010000110101111;
		correct = 32'b01110101110000001010000110101111;
		#400; //1.0731256e+22 * -4.8837907e+32 = 4.8837907e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001101011110110100100111000101;
		x2 = 32'b10111100100110111101001001000101;
		correct = 32'b00111100100110111101001001000101;
		#400; //7.7434143e-31 * -0.019021163 = 0.019021163
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011011100100010001111000010;
		x2 = 32'b10000010111000110100100101001000;
		correct = 32'b10000011000000000111111100011110;
		#400; //-7.1158456e-37 * -3.3396714e-37 = -3.7761743e-37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100101110010110000101101110;
		x2 = 32'b00011010001010000001100110001100;
		correct = 32'b11111100101110010110000101101110;
		#400; //-7.700408e+36 * 3.4762222e-23 = -7.700408e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011101001111011111101011000;
		x2 = 32'b10000010111111111110110111001100;
		correct = 32'b01001011101001111011111101011000;
		#400; //21986992.0 * -3.7605371e-37 = 21986992.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110110010010100011001101101110;
		x2 = 32'b11000011101001010110101001111011;
		correct = 32'b01000011101001010110101001111011;
		#400; //3.0130282e-06 * -330.83188 = 330.83188
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001000011100011101111010001000;
		x2 = 32'b00110001001110011011011110010010;
		correct = 32'b11001000011100011101111010001000;
		#400; //-247674.12 * 2.702539e-09 = -247674.12
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100100010100101100100111000;
		x2 = 32'b01111001100001110101001010111100;
		correct = 32'b11111001100001110101001010111100;
		#400; //-4753618600000.0 * 8.782977e+34 = -8.782977e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100110010101110011111101110;
		x2 = 32'b01001100000110000111111100001001;
		correct = 32'b11110100110010101110011111101110;
		#400; //-1.2860694e+32 * 39975972.0 = -1.2860694e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010001111110000111110110000111;
		x2 = 32'b10110000001001101111001011011100;
		correct = 32'b11010001111110000111110110000111;
		#400; //-133407240000.0 * -6.073557e-10 = -133407240000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011101100111100010110100101100;
		x2 = 32'b00100111100011100001001100011011;
		correct = 32'b01011101100111100010110100101100;
		#400; //1.4247268e+18 * 3.943363e-15 = 1.4247268e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100011111011101100010100100;
		x2 = 32'b01110100000000001101001101000010;
		correct = 32'b11111100011111011101100100100101;
		#400; //-5.2721804e+36 * 4.0826344e+31 = -5.2722213e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000110000000010001100101010;
		x2 = 32'b00110010000101101010100010000111;
		correct = 32'b11110000110000000010001100101010;
		#400; //-4.7570906e+29 * 8.769468e-09 = -4.7570906e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011011010101001111000111110100;
		x2 = 32'b11011010110110111001100000001000;
		correct = 32'b01011010110110111001100000001000;
		#400; //-1.7614408e-22 * -3.090509e+16 = 3.090509e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101101001110100001001101110011;
		x2 = 32'b01101101011111100001000001110111;
		correct = 32'b11101101110111000001000111110101;
		#400; //-3.5992328e+27 * 4.9143186e+27 = -8.5135514e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101101010010100100100010011;
		x2 = 32'b11111110111001011010001111010111;
		correct = 32'b01111110111001011010001111010111;
		#400; //0.08265891 * -1.5262196e+38 = 1.5262196e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100100111111011010011111011010;
		x2 = 32'b11100110110101111101011011011111;
		correct = 32'b01100110110001111111110001100001;
		#400; //-3.743297e+22 * -5.0963623e+23 = 4.7220325e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001111011101110011010001010011;
		x2 = 32'b00111110000100100001110100011110;
		correct = 32'b10111110000100100001110100011110;
		#400; //-1.21881175e-29 * 0.1426892 = -0.1426892
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101101100111111010110100110110;
		x2 = 32'b10011010111000001111110001001011;
		correct = 32'b01101101100111111010110100110110;
		#400; //6.1771895e+27 * -9.305183e-23 = 6.1771895e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101100001110000010001111001011;
		x2 = 32'b11101110000010001111010001100000;
		correct = 32'b01101101111110101110010001000111;
		#400; //-8.904455e+26 * -1.0596348e+28 = 9.705903e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010100000101100110111000111001;
		x2 = 32'b10100100100101000011100001100111;
		correct = 32'b01010100000101100110111000111001;
		#400; //2584377300000.0 * -6.428032e-17 = 2584377300000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000100010110010010111000011110;
		x2 = 32'b01011001110001011010100001001110;
		correct = 32'b11011001110001011010100001001110;
		#400; //-868.7206 * 6954453000000000.0 = -6954453000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000100111000100000100111111111;
		x2 = 32'b10011101101111101100110111000011;
		correct = 32'b00011101101111101100110111000011;
		#400; //5.3141525e-36 * -5.0505334e-21 = 5.0505334e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011101001001100111110100110;
		x2 = 32'b10100010111111111110011001100110;
		correct = 32'b01101011101001001100111110100110;
		#400; //3.9848885e+26 * -6.9361832e-18 = 3.9848885e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000011001101100101011010111010;
		x2 = 32'b01010101100001111111110111101001;
		correct = 32'b11010101100001111111110111101001;
		#400; //182.33878 * 18690576000000.0 = -18690576000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111001100000011011101001100100;
		x2 = 32'b11011000000101010100001011000010;
		correct = 32'b11111001100000011011101001100100;
		#400; //-8.419834e+34 * -656455800000000.0 = -8.419834e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101101001111111001100100110100;
		x2 = 32'b10100011100110110011101011010010;
		correct = 32'b00101101001111111001100101000111;
		#400; //1.0891111e-11 * -1.6830045e-17 = 1.0891127e-11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001100101101010010100110100011;
		x2 = 32'b11001010101011111011100100010111;
		correct = 32'b01001100110000000010010100110100;
		#400; //94981400.0 * -5758091.5 = 100739490.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101000101101101000001110010000;
		x2 = 32'b00011011001011001101101110110100;
		correct = 32'b11101000101101101000001110010000;
		#400; //-6.895181e+24 * 1.4298496e-22 = -6.895181e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000011100011000010001101111000;
		x2 = 32'b11011001111111111000111000101111;
		correct = 32'b01011001111111111000111000101111;
		#400; //8.236604e-37 * -8991556400000000.0 = 8991556400000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111111011111100000010000110111;
		x2 = 32'b10010101111011000110011111001000;
		correct = 32'b00111111011111100000010000110111;
		#400; //0.9922518 * -9.548338e-26 = 0.9922518
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010000110100001010001000011;
		x2 = 32'b00101110111101001111100011000000;
		correct = 32'b10101110111101010100010111001010;
		#400; //-1.3684977e-13 * 1.1140022e-10 = -1.1153707e-10
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111011011011010101010110011000;
		x2 = 32'b00001010110001110001111011000111;
		correct = 32'b10111011011011010101010110011000;
		#400; //-0.0036214348 * 1.917458e-32 = -0.0036214348
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011011111011100111111011101011;
		x2 = 32'b10110001111110111001101101100110;
		correct = 32'b00110001111110111001101101100110;
		#400; //3.9455816e-22 * -7.322728e-09 = 7.322728e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010011101001110100001110100111;
		x2 = 32'b00111110001011101011111011110000;
		correct = 32'b10111110001011101011111011110000;
		#400; //4.2223437e-27 * 0.17065024 = -0.17065024
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001001100011110101111000001;
		x2 = 32'b01010101100011110111101010001010;
		correct = 32'b11010101100011110111101010001010;
		#400; //3.950638e-14 * 19719558000000.0 = -19719558000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110001100011011100101100110011;
		x2 = 32'b01001110000000111001100001000101;
		correct = 32'b11110001100011011100101100110011;
		#400; //-1.4042573e+30 * 551948600.0 = -1.4042573e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101010001110010010110101000;
		x2 = 32'b10010101010110001001011010101000;
		correct = 32'b00110101010001110010010110101000;
		#400; //7.4188074e-07 * -4.37397e-26 = 7.4188074e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000110011010011101011111011001;
		x2 = 32'b11000100000001010110101000100101;
		correct = 32'b01000100000001010110101000100101;
		#400; //-4.398101e-35 * -533.6585 = 533.6585
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100011010010000000010011111;
		x2 = 32'b00011011100101111011010011001110;
		correct = 32'b10111100011010010000000010011111;
		#400; //-0.0142213395 * 2.5097697e-22 = -0.0142213395
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100010001011011001100110111;
		x2 = 32'b01100010111001000111111000101001;
		correct = 32'b01110100010001011011001100110111;
		#400; //6.265365e+31 * 2.1074742e+21 = 6.265365e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010000011110111001100011010010;
		x2 = 32'b11011111010100001011111010010111;
		correct = 32'b01011111010100001011111010010111;
		#400; //-4.961875e-29 * -1.5041626e+19 = 1.5041626e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100100001011011001011110011000;
		x2 = 32'b11111010100100011101100010101011;
		correct = 32'b01111010100100011101100010101011;
		#400; //-3.76418e-17 * -3.786388e+35 = 3.786388e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101111011100101111111100000;
		x2 = 32'b11010010111011011010001011011101;
		correct = 32'b01010010111011011010001011011101;
		#400; //0.116393805 * -510319820000.0 = 510319820000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000100100111000000011010011;
		x2 = 32'b00001100001000101101111111111110;
		correct = 32'b10011000100100111000000011010011;
		#400; //-3.812869e-24 * 1.2547431e-31 = -3.812869e-24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101111010110001101011100000000;
		x2 = 32'b01011010000011110011000010100111;
		correct = 32'b11011010000011110011000010100111;
		#400; //1.9721469e-10 * 1.0076104e+16 = -1.0076104e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011100000101000000110001011111;
		x2 = 32'b01000010100110000100000111000111;
		correct = 32'b11011100000101000000110001011111;
		#400; //-1.666876e+17 * 76.12847 = -1.666876e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100000101010110101101110011111;
		x2 = 32'b01101110010100110000010100100110;
		correct = 32'b11101110010100110000010100100110;
		#400; //2.9029157e-19 * 1.632689e+28 = -1.632689e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110000100001111011110100011;
		x2 = 32'b11001101110010010100010111101010;
		correct = 32'b01001101110010010100010111101010;
		#400; //-3.2961755e-11 * -422100300.0 = 422100300.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100001101101001100100000001;
		x2 = 32'b01110110101111110010100001101001;
		correct = 32'b11110110101111110010100001101001;
		#400; //-0.011144877 * 1.938571e+33 = -1.938571e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101000101011000000011101001;
		x2 = 32'b10001001010010101111101000110000;
		correct = 32'b11111101000101011000000011101001;
		#400; //-1.242027e+37 * -2.4432503e-33 = -1.242027e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111101101011011000000001101000;
		x2 = 32'b00111000010101110000000000000100;
		correct = 32'b10111101101011011001101101001000;
		#400; //-0.08471757 * 5.126001e-05 = -0.08476883
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000111101110000001101011001;
		x2 = 32'b01101111101111010101001110010000;
		correct = 32'b11110001000100110010110000011110;
		#400; //-6.1157476e+29 * 1.1718738e+29 = -7.287621e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111000001111111000011100111;
		x2 = 32'b00010010001101110010100000110111;
		correct = 32'b11111111000001111111000011100111;
		#400; //-1.8069662e+38 * 5.7794187e-28 = -1.8069662e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111000111011001110001001110001;
		x2 = 32'b01001100111010110111000100010001;
		correct = 32'b11001100111010110111000100010001;
		#400; //0.00011295535 * 123439240.0 = -123439240.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111010100100010001100011000001;
		x2 = 32'b11111000011010100101100100101101;
		correct = 32'b01111010100110000110101110001010;
		#400; //3.7669256e+35 * -1.9012596e+34 = 3.9570514e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001100011011100101001100011100;
		x2 = 32'b11000110000011110100011110000100;
		correct = 32'b01000110000011110100011110000100;
		#400; //-1.8359863e-31 * -9169.879 = 9169.879
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110110101011011011010111010010;
		x2 = 32'b11010101011010000101100000010111;
		correct = 32'b11110110101011011011010111010010;
		#400; //-1.761631e+33 * -15966565000000.0 = -1.761631e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000101101101001001000000001110;
		x2 = 32'b10101000011101001111011111000010;
		correct = 32'b11000101101101001001000000001110;
		#400; //-5778.007 * -1.3598445e-14 = -5778.007
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000111001001110111110011101001;
		x2 = 32'b00001000011101010011100010001110;
		correct = 32'b10001000100011111000101111100100;
		#400; //-1.2600391e-34 * 7.3793485e-34 = -8.639388e-34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100111010111010011100010010010;
		x2 = 32'b00101100111010110111101111111011;
		correct = 32'b11100111010111010011100010010010;
		#400; //-1.0446865e+24 * 6.6928663e-12 = -1.0446865e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111011101100001110101011101110;
		x2 = 32'b11001111010000011111111111110011;
		correct = 32'b01001111010000011111111111110011;
		#400; //0.0053990996 * -3254776600.0 = 3254776600.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000010110011110110111111011010;
		x2 = 32'b10110001111111101111100001001001;
		correct = 32'b00110001111111101111100001001001;
		#400; //-3.0480116e-37 * -7.4205997e-09 = 7.4205997e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100011110010101101000001011000;
		x2 = 32'b11111101100100110000100100001100;
		correct = 32'b01111101100100110000100100001100;
		#400; //-2.1989121e-17 * -2.4430436e+37 = 2.4430436e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111001011101100011010001010;
		x2 = 32'b11011110100100001110101111110000;
		correct = 32'b01011110100100001110101111110000;
		#400; //2.425498e-15 * -5.221352e+18 = 5.221352e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100100111010110101111100100;
		x2 = 32'b11011100111110100101011001100100;
		correct = 32'b01011100111110100101011001100100;
		#400; //-4.4741866e-12 * -5.6370985e+17 = 5.6370985e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000101111101111010100111011001;
		x2 = 32'b10111101100100000001011101010011;
		correct = 32'b01000101111101111010101001101001;
		#400; //7925.231 * -0.07035699 = 7925.3013
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001111000111100000100011110010;
		x2 = 32'b00100101000000000101000010100010;
		correct = 32'b01001111000111100000100011110010;
		#400; //2651386400.0 * 1.112955e-16 = 2651386400.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000100101001110111000110100110;
		x2 = 32'b01011111001001011010010001111110;
		correct = 32'b11011111001001011010010001111110;
		#400; //1339.5515 * 1.1935803e+19 = -1.1935803e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000100000010000010010000011111;
		x2 = 32'b11101001010010010011101101001101;
		correct = 32'b01101001010010010011101101001101;
		#400; //-544.5644 * -1.5204633e+25 = 1.5204633e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000110001011111011000100110;
		x2 = 32'b10101000001000000011100000010100;
		correct = 32'b00101000001000000011100000010100;
		#400; //7.808205e-29 * -8.893944e-15 = 8.893944e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011011111110000000100110000101;
		x2 = 32'b10011101001101010110101111011101;
		correct = 32'b00011101000101100110101010101100;
		#400; //-4.103431e-22 * -2.4010915e-21 = 1.9907483e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001001101010111110111001110001;
		x2 = 32'b00011010100001000101011110000110;
		correct = 32'b01001001101010111110111001110001;
		#400; //1408462.1 * 5.473532e-23 = 1408462.1
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101101000100010010111001101101;
		x2 = 32'b11011000101000000100011100000110;
		correct = 32'b01011000101000000100011100000110;
		#400; //8.252604e-12 * -1409815200000000.0 = 1409815200000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101101000111001111011010101;
		x2 = 32'b11101001000001001011000000001011;
		correct = 32'b01101001000001001011000000001011;
		#400; //0.07989279 * -1.0025597e+25 = 1.0025597e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110001101100100100101010000001;
		x2 = 32'b11110110011110001011101011111101;
		correct = 32'b01110110011110001011101011111101;
		#400; //5.188952e-09 * -1.2612131e+33 = 1.2612131e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001000000100011011001011000101;
		x2 = 32'b11110001011100111011111101010001;
		correct = 32'b01110001011100111011111101010001;
		#400; //4.3844493e-34 * -1.2069783e+30 = 1.2069783e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100010110110100110000010110001;
		x2 = 32'b00000001010011111110100111111111;
		correct = 32'b00100010110110100110000010110001;
		#400; //5.9191394e-18 * 3.818778e-38 = 5.9191394e-18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001100011000110100100101010001;
		x2 = 32'b11001101000010010100100101000010;
		correct = 32'b01001101000010010100100101000010;
		#400; //1.7509507e-31 * -143954980.0 = 143954980.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001011100110101110100100000101;
		x2 = 32'b00101101001110110010000111101100;
		correct = 32'b10101101001110110010000111101100;
		#400; //5.966925e-32 * 1.06372515e-11 = -1.06372515e-11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000010110111010001011010001111;
		x2 = 32'b11111100011100111111100111010000;
		correct = 32'b01111100011100111111100111010000;
		#400; //3.248598e-37 * -5.0671797e+36 = 5.0671797e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101011111000100100111111010011;
		x2 = 32'b01001010101100011110010000110111;
		correct = 32'b11001010101100011110010000110111;
		#400; //1.6080421e-12 * 5829147.5 = -5829147.5
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101111100001000000111100111001;
		x2 = 32'b00001010100111110010000010100010;
		correct = 32'b01101111100001000000111100111001;
		#400; //8.174085e+28 * 1.5323418e-32 = 8.174085e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101101110111010111110011111110;
		x2 = 32'b11101111010000100000110010011010;
		correct = 32'b01101111001001100101110011111010;
		#400; //-8.5684117e+27 * -6.0055326e+28 = 5.1486913e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110101101001001111101011000101;
		x2 = 32'b10001100001101100010000101010110;
		correct = 32'b11110101101001001111101011000101;
		#400; //-4.182729e+32 * -1.4030802e-31 = -4.182729e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101111101111111011010100000000;
		x2 = 32'b01011111001010001010110111010101;
		correct = 32'b01101111101111111011010100000000;
		#400; //1.18660905e+29 * 1.2154605e+19 = 1.18660905e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111000000101000101101111000101;
		x2 = 32'b10110010101001100110111101100010;
		correct = 32'b10111000000101000100011011110111;
		#400; //-3.5371417e-05 * -1.9375594e-08 = -3.535204e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110100011111011010010101111011;
		x2 = 32'b11110001000101011101100011010101;
		correct = 32'b01110001000101011101100011010101;
		#400; //-2.3622663e-07 * -7.420064e+29 = 7.420064e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100000011101010011010010101011;
		x2 = 32'b01010101011111110100011001000100;
		correct = 32'b01100000011101010011010010100111;
		#400; //7.067574e+19 * 17542328000000.0 = 7.0675723e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111001101010101011101101111;
		x2 = 32'b10110110100110011001001101010000;
		correct = 32'b11011111001101010101011101101111;
		#400; //-1.3067035e+19 * -4.5769048e-06 = -1.3067035e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000100010000010000110101111;
		x2 = 32'b01101010001010101100111101011010;
		correct = 32'b11101010001010101100111101011010;
		#400; //-3.5189188e-24 * 5.1624145e+25 = -5.1624145e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101101101001000010001100000010;
		x2 = 32'b10010100000000001111000000110010;
		correct = 32'b11101101101001000010001100000010;
		#400; //-6.349733e+27 * -6.509719e-27 = -6.349733e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111010000010011011001011110011;
		x2 = 32'b11100111001001110000111111110110;
		correct = 32'b11111010000010011011001011110011;
		#400; //-1.7874355e+35 * -7.889296e+23 = -1.7874355e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010010110001000111001110110100;
		x2 = 32'b01110111101100111111110011011010;
		correct = 32'b11110111101100111111110011011010;
		#400; //421877380000.0 * 7.3011686e+33 = -7.3011686e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000111110111111111001100101100;
		x2 = 32'b01010101100010101010010000000011;
		correct = 32'b11010101100010101010010000000011;
		#400; //-114662.34 * 19054629000000.0 = -19054629000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100001000110011101100110010;
		x2 = 32'b11101010011011111110111101000001;
		correct = 32'b01101010011011111110111101000001;
		#400; //-0.009962844 * -7.251578e+25 = 7.251578e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101011101010100100101111111;
		x2 = 32'b00011000011111001111001111101101;
		correct = 32'b10011000011111001111001111101101;
		#400; //1.1533344e-35 * 3.2693388e-24 = -3.2693388e-24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101101011100101101011101111001;
		x2 = 32'b10110110011001100110100111100001;
		correct = 32'b00110110011001100110100110100100;
		#400; //-1.3803952e-11 * -3.43343e-06 = 3.4334162e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100000100011010010101110100010;
		x2 = 32'b00110110100000001110111100101011;
		correct = 32'b10110110100000001110111100101011;
		#400; //-2.3915203e-19 * 3.84254e-06 = -3.84254e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110110000110011110110100101010;
		x2 = 32'b01110111011010011011001011101001;
		correct = 32'b11110111011010011011001011101001;
		#400; //2.2936824e-06 * 4.7399762e+33 = -4.7399762e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000000110111101001010101101010;
		x2 = 32'b11011000001010110100100101101111;
		correct = 32'b01011000001010110100100101101111;
		#400; //-2.044108e-38 * -753327500000000.0 = 753327500000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001000110010001111101111001110;
		x2 = 32'b11100101000010001111101100001110;
		correct = 32'b01100101000010001111101100001110;
		#400; //1.2096261e-33 * -4.042956e+22 = 4.042956e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010010100011101000100000010;
		x2 = 32'b00100001110111100011000101101110;
		correct = 32'b10101010010100011101000101110001;
		#400; //-1.8635443e-13 * 1.5056389e-18 = -1.8635594e-13
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001110111011110101011000111000;
		x2 = 32'b01110011010100101111110011111000;
		correct = 32'b11110011010100101111110011111000;
		#400; //5.9001074e-30 * 1.6716204e+31 = -1.6716204e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100111101011011110101110000101;
		x2 = 32'b01100010000100000001111010110010;
		correct = 32'b11100010000100000001111010110010;
		#400; //-4.8272497e-15 * 6.6463574e+20 = -6.6463574e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101101000000000110101011111101;
		x2 = 32'b10101100001100111110100001100110;
		correct = 32'b00101101001011010110010100010110;
		#400; //7.299714e-12 * -2.5566437e-12 = 9.856357e-12
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011100010101101101001110101001;
		x2 = 32'b00101000111110100111110100001110;
		correct = 32'b10101000111110100111110100001110;
		#400; //7.1080225e-22 * 2.780981e-14 = -2.780981e-14
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000000101011011100000110000110;
		x2 = 32'b10101111100000000010000111110101;
		correct = 32'b01000000101011011100000110000110;
		#400; //5.4298735 * -2.3307192e-10 = 5.4298735
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000100100101111011010111101000;
		x2 = 32'b00101001100111111100001100001110;
		correct = 32'b10101001100111111100001100001110;
		#400; //-3.5666984e-36 * 7.094855e-14 = -7.094855e-14
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110010100011000110001101101110;
		x2 = 32'b00110111000010101000100000101001;
		correct = 32'b11110010100011000110001101101110;
		#400; //-5.5613574e+30 * 8.257143e-06 = -5.5613574e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101100100101011001010000010001;
		x2 = 32'b11001110000100101001110000000011;
		correct = 32'b01001110000100101001110000000011;
		#400; //4.2512734e-12 * -614924500.0 = 614924500.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100111101101000110010000101110;
		x2 = 32'b11011101011001001001101110010010;
		correct = 32'b01011101011001001001101110010010;
		#400; //-5.006865e-15 * -1.02955754e+18 = 1.02955754e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110001111011000110100001011111;
		x2 = 32'b01011101101111000101110000100111;
		correct = 32'b11011101101111000101110000100111;
		#400; //6.8803696e-09 * 1.6965958e+18 = -1.6965958e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111001010110111101100011100011;
		x2 = 32'b11010001111001100000001101111101;
		correct = 32'b01010001111001100000001101111101;
		#400; //0.00020966264 * -123487625000.0 = 123487625000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101110000010100101100101011110;
		x2 = 32'b11001010000001111000010000110111;
		correct = 32'b01101110000010100101100101011110;
		#400; //1.0704242e+28 * -2220301.8 = 1.0704242e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101101110101010011101100011;
		x2 = 32'b00100101010101000110001010111111;
		correct = 32'b00111101101110101010011101100011;
		#400; //0.09113958 * 1.8421525e-16 = 0.09113958
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101110110111110001110000000100;
		x2 = 32'b01100000011100101111100100110000;
		correct = 32'b11101110110111110001110000000100;
		#400; //-3.4524513e+28 * 7.003231e+19 = -3.4524513e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101010011110101010001111101;
		x2 = 32'b11100111011100000001101110011001;
		correct = 32'b01100111011100000001101110011001;
		#400; //-1.7983014e-16 * -1.13387704e+24 = 1.13387704e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000011100110111011000001111000;
		x2 = 32'b01000101000001100100000011011000;
		correct = 32'b11000101000001100100000011011000;
		#400; //9.1505965e-37 * 2148.0527 = -2148.0527
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001110100111101111001011010011;
		x2 = 32'b10000010101000111101110110010000;
		correct = 32'b01001110100111101111001011010011;
		#400; //1333356900.0 * -2.4077868e-37 = 1333356900.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000110101001000111010111110101;
		x2 = 32'b11100001111011101000011001110101;
		correct = 32'b01100001111011101000011001110101;
		#400; //21050.979 * -5.500017e+20 = 5.500017e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110111011000011001111000111;
		x2 = 32'b01101000001100101011011110100100;
		correct = 32'b11101000001100101011011110100100;
		#400; //8.8849413e-35 * 3.3758752e+24 = -3.3758752e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100100001101001100101001010101;
		x2 = 32'b11101001010110110101010100000110;
		correct = 32'b01101001010110110101010100000110;
		#400; //-3.920266e-17 * -1.6572267e+25 = 1.6572267e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100000100001000100000111110000;
		x2 = 32'b01001110001011001100110011000110;
		correct = 32'b11001110001011001100110011000110;
		#400; //-2.2405304e-19 * 724775300.0 = -724775300.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101100110001010010111101000;
		x2 = 32'b11001110000111000011101010000001;
		correct = 32'b11111101100110001010010111101000;
		#400; //-2.536301e+37 * -655269950.0 = -2.536301e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110111000001000111011010110;
		x2 = 32'b01101110001111110100010001110010;
		correct = 32'b11101110001111110100010001110010;
		#400; //-1.02117134e-10 * 1.4798596e+28 = -1.4798596e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101110100100101001010100111101;
		x2 = 32'b00111100001011010001000111011110;
		correct = 32'b10111100001011010001000111011110;
		#400; //6.6658214e-11 * 0.010563342 = -0.010563342
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010100100011011110011000100110;
		x2 = 32'b10011110100010011101111001000001;
		correct = 32'b01010100100011011110011000100110;
		#400; //4875613000000.0 * -1.4597361e-20 = 4875613000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001101101001000000110100100000;
		x2 = 32'b10111100110111000110100011110110;
		correct = 32'b00111100110111000110100011110110;
		#400; //1.011044e-30 * -0.026905518 = 0.026905518
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010100110000101001010100011;
		x2 = 32'b10000111100100110011110110010001;
		correct = 32'b01000010100110000101001010100011;
		#400; //76.1614 * -2.2154287e-34 = 76.1614
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111010001101111000110011110;
		x2 = 32'b10101011100011000001010000010101;
		correct = 32'b11010111010001101111000110011110;
		#400; //-218741040000000.0 * -9.953172e-13 = -218741040000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000100101110110010111110111000;
		x2 = 32'b11001010011111000111100010101110;
		correct = 32'b01001010011111000110000101001000;
		#400; //-1497.4912 * -4136491.5 = 4134994.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000101011110111111110100100100;
		x2 = 32'b10011100001100001110000110010011;
		correct = 32'b00011100001100001110000110010011;
		#400; //-1.1848458e-35 * -5.8525063e-22 = 5.8525063e-22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000101101001010110111000111111;
		x2 = 32'b00111001010011010110110000101011;
		correct = 32'b01000101101001010110111000111111;
		#400; //5293.781 * 0.00019590619 = 5293.781
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111000100100010100111011100011;
		x2 = 32'b00010010111110011001111111101110;
		correct = 32'b10111000100100010100111011100011;
		#400; //-6.9288326e-05 * 1.5753535e-27 = -6.9288326e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110010100111111000101001010101;
		x2 = 32'b10011011000100111011110110011010;
		correct = 32'b01110010100111111000101001010101;
		#400; //6.320045e+30 * -1.2220819e-22 = 6.320045e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011110011001110011101110110111;
		x2 = 32'b01011111100101111110000000100111;
		correct = 32'b11011111100101111110000000100111;
		#400; //1.2241387e-20 * 2.188758e+19 = -2.188758e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111010000011010011100100000100;
		x2 = 32'b01001011001001001101000000000111;
		correct = 32'b11001011001001001101000000000111;
		#400; //-0.0005387219 * 10801159.0 = -10801159.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011111101100101101100101011;
		x2 = 32'b11111001100110011110010110011010;
		correct = 32'b01111001100110011110010110011010;
		#400; //-1.4479512e-36 * -9.988479e+34 = 9.988479e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110000100111000110110110011;
		x2 = 32'b01000011100001010001101100110001;
		correct = 32'b11000011100001010000100010111111;
		#400; //0.14409523 * 266.21243 = -266.06833
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010011000100010111111111011101;
		x2 = 32'b00111110110111000101110001101001;
		correct = 32'b10111110110111000101110001101001;
		#400; //-1.8364614e-27 * 0.43039253 = -0.43039253
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001011001111101011011110111010;
		x2 = 32'b01000000101000100001000010100110;
		correct = 32'b11001011001111101011011110111111;
		#400; //-12498874.0 * 5.0645323 = -12498879.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100010101000010101011111111000;
		x2 = 32'b10111101100100101110111010000110;
		correct = 32'b00111101100100101110111010000110;
		#400; //4.373228e-18 * -0.07174401 = 0.07174401
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110111000101000101000111000110;
		x2 = 32'b11100110010000110111111111011110;
		correct = 32'b01110111000101000101000111000110;
		#400; //3.0082754e+33 * -2.3080505e+23 = 3.0082754e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100010011110111111011100001010;
		x2 = 32'b10000001000001011000000001111000;
		correct = 32'b11100010011110111111011100001010;
		#400; //-1.16198345e+21 * -2.4520414e-38 = -1.16198345e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111001010111111100011000001110;
		x2 = 32'b10010011100001101111111000001111;
		correct = 32'b11111001010111111100011000001110;
		#400; //-7.26187e+34 * -3.4076877e-27 = -7.26187e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end
end
endmodule