`timescale 1 ns/1 ps
    `include "alu.v"


    module add_tb ();
        reg clk;
        reg [31:0] x1, x2;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] x3;
        wire [49:0] pro;

        alu U1 (
                .clk(clk),
                .x1(x1),
                .x2(x2),
                .OpCode(op),
                .x3(x3)
            );
        
        always
        #200 clk = ~clk; 
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clk, x1, x2, op, x3);
            clk = 0;

    op = 3'b000;

		
		$display ("Opcode -> 000, Operation -> ADD");
		
		
		x1 = 32'b10110111001001011010001101000111;
		x2 = 32'b01000111110110100100000110001001;
		correct = 32'b01000111110110100100000110001001;
		#500; //-9.872782e-06 * 111747.07 = 111747.07
					begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001101110110101101010101101001;
		x2 = 32'b01011010010101101100100000000000;
		correct = 32'b01011010010101101100100000000000;
		#500; //458927400.0 * 1.5113887e+16 = 1.5113887e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001110000100111100111101100;
		x2 = 32'b10011011001001011111100001111001;
		correct = 32'b11000001110000100111100111101100;
		#500; //-24.309532 * -1.3728766e-22 = -24.309532
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101111110001111000010111010;
		x2 = 32'b00011000000011100000110011100101;
		correct = 32'b00110101111110001111000010111010;
		#500; //1.85475e-06 * 1.835958e-24 = 1.85475e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100010110010111011101101111110;
		x2 = 32'b11101010101010011100110101011100;
		correct = 32'b11101010101010011100111000101000;
		#500; //-1.8790996e+21 * -1.0263912e+26 = -1.02641e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001000110011000110000011101000;
		x2 = 32'b01010011000011001010110010000010;
		correct = 32'b01010011000011001010110010001000;
		#500; //418567.25 * 604189600000.0 = 604190000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100111000000110110010010011;
		x2 = 32'b10101001101111000000001000100101;
		correct = 32'b00111100111000000110110010010011;
		#500; //0.027395522 * -8.349249e-14 = 0.027395522
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011001001101101111001110100;
		x2 = 32'b01111011101110011100000011101010;
		correct = 32'b01111011101110011100000011101010;
		#500; //2.017322e+26 * 1.9289754e+36 = 1.9289754e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101101100111000100111010000;
		x2 = 32'b10100010001000001111111011100100;
		correct = 32'b00110101101100111000100111010000;
		#500; //1.3376648e-06 * -2.1818981e-18 = 1.3376648e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010101011110010010101101110011;
		x2 = 32'b10000110100000001001100110101001;
		correct = 32'b10010101011110010010101101110011;
		#500; //-5.0319425e-26 * -4.837403e-35 = -5.0319425e-26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100000011100001011000100011;
		x2 = 32'b10111010001101110011010001101100;
		correct = 32'b10111100000110011000100101101010;
		#500; //-0.00867227 * -0.00069887075 = -0.009371141
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010110111000100001111001111101;
		x2 = 32'b01010001011111001010000011000100;
		correct = 32'b01010001011111001010000011000100;
		#500; //3.653151e-25 * 67814310000.0 = 67814310000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100000110101100101111100000;
		x2 = 32'b01110100000110111000111101111010;
		correct = 32'b01110100000110111000111101111010;
		#500; //-5.121783e-22 * 4.9299076e+31 = 4.9299076e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001100010100001100011010111101;
		x2 = 32'b00110110101110010111000101011111;
		correct = 32'b01001100010100001100011010111101;
		#500; //54729460.0 * 5.526628e-06 = 54729460.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101011100101110111101100010000;
		x2 = 32'b00000111000010110100110110101011;
		correct = 32'b11101011100101110111101100010000;
		#500; //-3.662579e+26 * 1.0480022e-34 = -3.662579e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000010011111001010001110110110;
		x2 = 32'b01111101100011100111111011011000;
		correct = 32'b01111101100011100111111011011000;
		#500; //-63.159874 * 2.3676123e+37 = 2.3676123e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010110000011100101011000101011;
		x2 = 32'b00001010011100000110011011000100;
		correct = 32'b11010110000011100101011000101011;
		#500; //-39125185000000.0 * 1.1574908e-32 = -39125185000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010010110011000111011111101101;
		x2 = 32'b10000011001000100101000100001100;
		correct = 32'b01010010110011000111011111101101;
		#500; //439092670000.0 * -4.770056e-37 = 439092670000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101010111011101010101111011101;
		x2 = 32'b11001011011011111011111110001010;
		correct = 32'b11101010111011101010101111011101;
		#500; //-1.4426797e+26 * -15712138.0 = -1.4426797e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110101100101000000101110111;
		x2 = 32'b11000010101001001011110011100111;
		correct = 32'b11111110101100101000000101110111;
		#500; //-1.186374e+38 * -82.36895 = -1.186374e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110110000010000010000101011011;
		x2 = 32'b10001001011000100111011001000110;
		correct = 32'b11110110000010000010000101011011;
		#500; //-6.902626e+32 * -2.7259372e-33 = -6.902626e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101010000011010010010100011111;
		x2 = 32'b00010111111101101011001101110000;
		correct = 32'b01101010000011010010010100011111;
		#500; //4.265846e+25 * 1.5942674e-24 = 4.265846e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010011011111111110010010010101;
		x2 = 32'b11000111001001011111010001110011;
		correct = 32'b11000111001001011111010001110011;
		#500; //-3.2298225e-27 * -42484.45 = -42484.45
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011011111111001001011101101101;
		x2 = 32'b00010010101000000000110010000000;
		correct = 32'b00011011111111001001011110010101;
		#500; //4.178776e-22 * 1.0100501e-27 = 4.178786e-22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001011011011111000001101001001;
		x2 = 32'b00110010100111100101000101101001;
		correct = 32'b00110010100111100101000101101001;
		#500; //-4.6128494e-32 * 1.8430642e-08 = 1.8430642e-08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101111010101001100001000110;
		x2 = 32'b11101001011100000000011010100001;
		correct = 32'b01111101111010101001100001000110;
		#500; //3.897875e+37 * -1.8135844e+25 = 3.897875e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110111101100111001010111110111;
		x2 = 32'b00100111100001000110110110111001;
		correct = 32'b11110111101100111001010111110111;
		#500; //-7.2848655e+33 * 3.675632e-15 = -7.2848655e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010011101100010010010000110111;
		x2 = 32'b00011100101111110100111110110110;
		correct = 32'b01010011101100010010010000110111;
		#500; //1521633600000.0 * 1.2659925e-21 = 1521633600000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011011101101111010000100111110;
		x2 = 32'b00011011100000111010111111000000;
		correct = 32'b10011010110011111100010111111000;
		#500; //-3.037901e-22 * 2.1785708e-22 = -8.593303e-23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001111101100100001001001010;
		x2 = 32'b00000110001000010101100000111001;
		correct = 32'b01111001111101100100001001001010;
		#500; //1.5983119e+35 * 3.034555e-35 = 1.5983119e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011011111101010010001001011000;
		x2 = 32'b10010010000010000101101110111010;
		correct = 32'b00011011111101010010001001000111;
		#500; //4.0554044e-22 * -4.3027095e-28 = 4.0554e-22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101111110010101110101000010;
		x2 = 32'b00101001001111001100101101110111;
		correct = 32'b00101001001111001100101101110111;
		#500; //2.3450105e-35 * 4.1920863e-14 = 4.1920863e-14
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100011101000100010001111111;
		x2 = 32'b11110111000001011010100100010011;
		correct = 32'b11110111000001011010100100010011;
		#500; //0.014908909 * -2.710956e+33 = -2.710956e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110000110010011111101011011000;
		x2 = 32'b01010010001110100011100010001101;
		correct = 32'b01010010001110100011100010001101;
		#500; //-1.4695969e-09 * 199953170000.0 = 199953170000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111100011000110101001010001111;
		x2 = 32'b00011001011101110001101110100101;
		correct = 32'b01111100011000110101001010001111;
		#500; //4.7213035e+36 * 1.27751835e-23 = 4.7213035e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001110001101100000101100110001;
		x2 = 32'b10111011110001000101110100011001;
		correct = 32'b01001110001101100000101100110001;
		#500; //763546700.0 * -0.0059925434 = 763546700.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011001000111001111011111010101;
		x2 = 32'b00100110101010100101011111010010;
		correct = 32'b11011001000111001111011111010101;
		#500; //-2761412000000000.0 * 1.1819923e-15 = -2761412000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011111101100101011111111101001;
		x2 = 32'b11001000110101100011011011010101;
		correct = 32'b11001000110101100011011011010101;
		#500; //7.570342e-20 * -438710.66 = -438710.66
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110010110011010111110101100010;
		x2 = 32'b00010110111011000101000111100101;
		correct = 32'b10110010110011010111110101100010;
		#500; //-2.3922158e-08 * 3.817954e-25 = -2.3922158e-08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000011111101101010101011001011;
		x2 = 32'b11000101100110110100000011000111;
		correct = 32'b11000101100010111101011000011010;
		#500; //493.33432 * -4968.097 = -4474.7627
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001110011010101000011101001001;
		x2 = 32'b00110110010111100101100101111111;
		correct = 32'b00110110010111100101100101111111;
		#500; //2.8907864e-30 * 3.3132671e-06 = 3.3132671e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110010111101111000101101001001;
		x2 = 32'b00100000000110111001010101111100;
		correct = 32'b01110010111101111000101101001001;
		#500; //9.8062314e+30 * 1.3178471e-19 = 9.8062314e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011011100110101111101010010;
		x2 = 32'b10100110110111110101110100111111;
		correct = 32'b10100110110111110101110100111111;
		#500; //-7.1520704e-37 * -1.5499008e-15 = -1.5499008e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000000010000000011100100010101;
		x2 = 32'b00110101100100010000111110011111;
		correct = 32'b11000000010000000011100100010000;
		#500; //-3.003484 * 1.0807888e-06 = -3.0034828
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001000111001001000010011100000;
		x2 = 32'b10100110001110111011001100111010;
		correct = 32'b10100110001110111011001100111010;
		#500; //-1.375349e-33 * -6.5121555e-16 = -6.5121555e-16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100101000111010101100100000100;
		x2 = 32'b10010101111110000000110111111111;
		correct = 32'b11100101000111010101100100000100;
		#500; //-4.644085e+22 * -1.00188484e-25 = -4.644085e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000100010001110111100100011;
		x2 = 32'b11010010111110110001010101001110;
		correct = 32'b11110000100010001110111100100011;
		#500; //-3.3903248e+29 * -539197100000.0 = -3.3903248e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000101010100000000001101001001;
		x2 = 32'b01001000010010010100011101001100;
		correct = 32'b01001000010010010100011101001100;
		#500; //-9.7807164e-36 * 206109.19 = 206109.19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101110000000010010101001101100;
		x2 = 32'b11010000000001111100001010111000;
		correct = 32'b11010000000001111100001010111000;
		#500; //2.9368882e-11 * -9110741000.0 = -9110741000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011101010111000001011101100;
		x2 = 32'b10111111011101000101010010000101;
		correct = 32'b10111111011101000101010010000101;
		#500; //1.8595305e-17 * -0.95441467 = -0.95441467
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100010011110111101011101100110;
		x2 = 32'b11100001101101111010100001001100;
		correct = 32'b11100001101101111010100001001100;
		#500; //3.4130874e-18 * -4.2348515e+20 = -4.2348515e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011111010110010101001101000110;
		x2 = 32'b01011110000111100001010000010001;
		correct = 32'b01011111100000000110110000100101;
		#500; //1.5659937e+19 * 2.847687e+18 = 1.8507624e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001000111100000010100010001111;
		x2 = 32'b10111011101001001011110101001100;
		correct = 32'b10111011101001001011110101001100;
		#500; //1.445401e-33 * -0.0050274488 = -0.0050274488
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100101010110111110011111000011;
		x2 = 32'b01101100001101001011111010111011;
		correct = 32'b01101100001101001011101101001011;
		#500; //-6.4904594e+22 * 8.740294e+26 = 8.7396445e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111100110000110011100100111;
		x2 = 32'b11011011110101011100110111000011;
		correct = 32'b11011011110101011100110111000011;
		#500; //1.8167846e-05 * -1.20360815e+17 = -1.20360815e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100100010111100000001101011;
		x2 = 32'b11100110110111101111110011001100;
		correct = 32'b01110100100010111100000001101011;
		#500; //8.857812e+31 * -5.2651432e+23 = 8.857812e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111001001100111111110100101000;
		x2 = 32'b00010000000000001001100101001011;
		correct = 32'b11111001001100111111110100101000;
		#500; //-5.8409735e+34 * 2.5361642e-29 = -5.8409735e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000110011111101101010000100;
		x2 = 32'b01101110111010011011100011100000;
		correct = 32'b11110000110000010011111011110110;
		#500; //-5.1462053e+29 * 3.6166754e+28 = -4.7845378e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011000101011011011001100111;
		x2 = 32'b11011010011001101000011000011011;
		correct = 32'b11111011000101011011011001100111;
		#500; //-7.773518e+35 * -1.6221674e+16 = -7.773518e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010001100001100110010101001010;
		x2 = 32'b01011000011110010111011001100101;
		correct = 32'b01011000011110010111001000110010;
		#500; //-72153120000.0 * 1097147600000000.0 = 1097075440000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011011000011001100100011000100;
		x2 = 32'b00111100011001111000011011001000;
		correct = 32'b01011011000011001100100011000100;
		#500; //3.962724e+16 * 0.014131255 = 3.962724e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100001100011110101100000111;
		x2 = 32'b00001101011110100001111101001110;
		correct = 32'b10111100001100011110101100000111;
		#500; //-0.010859258 * 7.707488e-31 = -0.010859258
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111011110101010110100001101010;
		x2 = 32'b10100011110110111111110111000011;
		correct = 32'b00111011110101010110100001101010;
		#500; //0.0065126913 * -2.38515e-17 = 0.0065126913
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111100001011111100010110010;
		x2 = 32'b11001010101101000101001101100101;
		correct = 32'b11001010101101000101001101100101;
		#500; //3.718455e-15 * -5908914.5 = -5908914.5
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001000101001111110011101111110;
		x2 = 32'b11010001100010100001000110101010;
		correct = 32'b11010001100010100001000110000000;
		#500; //343867.94 * -74125230000.0 = -74124890000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110000011010110011000101101110;
		x2 = 32'b10000101101101101111011100111100;
		correct = 32'b00110000011010110011000101101110;
		#500; //8.5562746e-10 * -1.7206017e-35 = 8.5562746e-10
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001000000101011000100010000001;
		x2 = 32'b11100101100101010110111011111111;
		correct = 32'b11100101100101010110111011111111;
		#500; //-153122.02 * -8.8210015e+22 = -8.8210015e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100011000110010111010010110111;
		x2 = 32'b10011010011010011100010000111101;
		correct = 32'b11100011000110010111010010110111;
		#500; //-2.830762e+21 * -4.834179e-23 = -2.830762e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000010000000101110100101110000;
		x2 = 32'b01011100110010111011000011100001;
		correct = 32'b01011100110010111011000011100001;
		#500; //9.617885e-38 * 4.586712e+17 = 4.586712e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101110000100111110001111101110;
		x2 = 32'b00000000110000001011111100111111;
		correct = 32'b01101110000100111110001111101110;
		#500; //1.1442462e+28 * 1.7701021e-38 = 1.1442462e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100100110100000101011001111111;
		x2 = 32'b11010100010000010000101101001011;
		correct = 32'b01100100110100000101011001111111;
		#500; //3.0745244e+22 * -3316472600000.0 = 3.0745244e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010000111101110111011110000100;
		x2 = 32'b10000101110011000001101110000110;
		correct = 32'b11010000111101110111011110000100;
		#500; //-33214440000.0 * -1.9194178e-35 = -33214440000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100111001101011100011000001100;
		x2 = 32'b01000101101111111000111010010110;
		correct = 32'b01100111001101011100011000001100;
		#500; //8.5840165e+23 * 6129.823 = 8.5840165e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010111111100101000000000001110;
		x2 = 32'b00100001001000110011011011110100;
		correct = 32'b00100001001000110011011100010010;
		#500; //1.5671209e-24 * 5.529928e-19 = 5.5299433e-19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101010111010011111110010000;
		x2 = 32'b11001100100010101110110010110101;
		correct = 32'b11001100100010101110110010110101;
		#500; //0.054015696 * -72836520.0 = -72836520.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110101011011011010111000010;
		x2 = 32'b00111001100011011101111010011101;
		correct = 32'b00111001100011011101111010011010;
		#500; //-7.899416e-11 * 0.00027059476 = 0.00027059467
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001001101000100001001010001110;
		x2 = 32'b01010001000101000111011001111010;
		correct = 32'b01010001000101000111011001111010;
		#500; //3.901753e-33 * 39852680000.0 = 39852680000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100111000111100001100000000000;
		x2 = 32'b10010111011001111111010101100000;
		correct = 32'b10100111000111100001100000000000;
		#500; //-2.1939915e-15 * -7.494983e-25 = -2.1939915e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010010001000101100011111011100;
		x2 = 32'b11000101000101101110010011010000;
		correct = 32'b11000101000101101110010011010000;
		#500; //-5.136453e-28 * -2414.3008 = -2414.3008
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000010011011111111110100100011;
		x2 = 32'b11001101010010010101001101001110;
		correct = 32'b11001101010010010101001101010010;
		#500; //-59.997204 * -211105000.0 = -211105060.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000110100000110111101011001010;
		x2 = 32'b11001110111100011100010101100100;
		correct = 32'b11001110111100011100010011100001;
		#500; //16829.395 * -2028122600.0 = -2028105900.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011000111100011001101011111010;
		x2 = 32'b10001010011010111101011011100110;
		correct = 32'b11011000111100011001101011111010;
		#500; //-2125183400000000.0 * -1.1355256e-32 = -2125183400000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101010000010011011100110100101;
		x2 = 32'b00001110010101000010000101111101;
		correct = 32'b00101010000010011011100110100101;
		#500; //1.2232453e-13 * 2.6147142e-30 = 1.2232453e-13
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110000101101110110001110110;
		x2 = 32'b00100011110110010110001100010011;
		correct = 32'b00100011110110010110001100010011;
		#500; //2.8385588e-35 * 2.3569147e-17 = 2.3569147e-17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011110010010111000110101011110;
		x2 = 32'b00001001111000001000000010000001;
		correct = 32'b01011110010010111000110101011110;
		#500; //3.6668707e+18 * 5.4046883e-33 = 3.6668707e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100011111111110100011111000110;
		x2 = 32'b10011111110101110010110001101100;
		correct = 32'b01100011111111110100011111000110;
		#500; //9.418183e+21 * -9.112953e-20 = 9.418183e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100101100100000000000000101011;
		x2 = 32'b01100000011011000001010111101000;
		correct = 32'b01100000011011000001010111101000;
		#500; //2.4980132e-16 * 6.8047033e+19 = 6.8047033e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101010001000000010000001100000;
		x2 = 32'b10100000000010000110101110011001;
		correct = 32'b11101010001000000010000001100000;
		#500; //-4.8395254e+25 * -1.1555249e-19 = -4.8395254e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101110100001111110010000111;
		x2 = 32'b01011010001111100110010110001110;
		correct = 32'b01110101110100001111110010000111;
		#500; //5.2984356e+32 * 1.3397977e+16 = 5.2984356e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000111010111100101111111111110;
		x2 = 32'b01010010111110110011011001101100;
		correct = 32'b01010010111110110011011001101100;
		#500; //-1.6729633e-34 * 539474920000.0 = 539474920000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011111001100101001011100011000;
		x2 = 32'b11010000111110010000101001010011;
		correct = 32'b11010000111110010000101001010011;
		#500; //3.7817948e-20 * -33425627000.0 = -33425627000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000111110000010110110110011010;
		x2 = 32'b10101000100010111010111000011111;
		correct = 32'b10101000100010111010111000011111;
		#500; //2.910383e-34 * -1.5507613e-14 = -1.5507613e-14
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110010001101110010000111000001;
		x2 = 32'b10000001100000010101011111010011;
		correct = 32'b10110010001101110010000111000001;
		#500; //-1.0659677e-08 * -4.751314e-38 = -1.0659677e-08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100011100000100101001011011;
		x2 = 32'b11011010110111111100101110100110;
		correct = 32'b01110100011100000100101001011011;
		#500; //7.6151084e+31 * -3.1496417e+16 = 7.6151084e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101000010010000000111101110;
		x2 = 32'b00100101010011011100011110100101;
		correct = 32'b01110101000010010000000111101110;
		#500; //1.7367769e+32 * 1.7848558e-16 = 1.7367769e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001111000010001111111110111110;
		x2 = 32'b11001011100100000100010010100101;
		correct = 32'b11001011100100000100010010100101;
		#500; //-6.754572e-30 * -18909514.0 = -18909514.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111100100000001100000101100001;
		x2 = 32'b11111111001111001001100111110010;
		correct = 32'b11111111001110001001001111100111;
		#500; //5.3482895e+36 * -2.506942e+38 = -2.453459e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110010011110010111100011011011;
		x2 = 32'b11100010010110010110011101010110;
		correct = 32'b11100010010110010110011101010110;
		#500; //-1.4521187e-08 * -1.0025974e+21 = -1.0025974e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001100100101001101101100110010;
		x2 = 32'b00101011011101100001111100111011;
		correct = 32'b00101011011101100001111100111011;
		#500; //2.2934934e-31 * 8.74401e-13 = 8.74401e-13
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111010011000101110101000000010;
		x2 = 32'b01000110110001100110110101110100;
		correct = 32'b11111010011000101110101000000010;
		#500; //-2.9455133e+35 * 25398.727 = -2.9455133e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111010010011011101110000010100;
		x2 = 32'b00011010110110111001111001000001;
		correct = 32'b10111010010011011101110000010100;
		#500; //-0.00078529236 * 9.083195e-23 = -0.00078529236
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100110000010101110100110011;
		x2 = 32'b11000011011001110011100000010010;
		correct = 32'b11000011011001110011100000010010;
		#500; //-1.952478e-26 * -231.21902 = -231.21902
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110100110100101001000110010;
		x2 = 32'b11110110110100101110001011010000;
		correct = 32'b11110110110100101110001011010000;
		#500; //5.8049137e-35 * -2.138638e+33 = -2.138638e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100010000101000001000111011001;
		x2 = 32'b10010010001111101111010101011000;
		correct = 32'b00100010000101000001000111011001;
		#500; //2.0067189e-18 * -6.025584e-28 = 2.0067189e-18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010110000111111000111111010101;
		x2 = 32'b01110110010100001111010011011010;
		correct = 32'b01110110010100001111010011011010;
		#500; //-1.2889303e-25 * 1.0595351e+33 = 1.0595351e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000100010010101001111001001101;
		x2 = 32'b00001010010000001100010010101000;
		correct = 32'b11000100010010101001111001001101;
		#500; //-810.47345 * 9.281451e-33 = -810.47345
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101000011000110000100111111;
		x2 = 32'b00111101101011001001100011001101;
		correct = 32'b11111101000011000110000100111111;
		#500; //-1.1662303e+37 * 0.08427582 = -1.1662303e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100010000111010010000000100111;
		x2 = 32'b11110100110010111000101100101011;
		correct = 32'b11110100110010111000101100101011;
		#500; //-7.246139e+20 * -1.290111e+32 = -1.290111e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101011111110100100110111100111;
		x2 = 32'b00001000000010100011110101111000;
		correct = 32'b11101011111110100100110111100111;
		#500; //-6.0519868e+26 * 4.160012e-34 = -6.0519868e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100001011000100101110000100111;
		x2 = 32'b00101010100101100001001111010101;
		correct = 32'b01100001011000100101110000100111;
		#500; //2.6097528e+20 * 2.6659114e-13 = 2.6097528e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000111010000010111110100111011;
		x2 = 32'b00010010011001010010111000110111;
		correct = 32'b11000111010000010111110100111011;
		#500; //-49533.23 * 7.2316623e-28 = -49533.23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000111000011011101100110111;
		x2 = 32'b00011110000110100101000010111011;
		correct = 32'b00011110000110100011010010000100;
		#500; //-5.8350176e-24 * 8.169387e-21 = 8.163552e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001111001000011001110001100111;
		x2 = 32'b01001000100111000110110100100111;
		correct = 32'b11001111001000011001011110000100;
		#500; //-2711381800.0 * 320361.22 = -2711061500.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111010011001010101001111111011;
		x2 = 32'b00100100101011011111110111110110;
		correct = 32'b10111010011001010101001111111011;
		#500; //-0.0008748171 * 7.545702e-17 = -0.0008748171
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000011111011001011111110011100;
		x2 = 32'b11100101111100010011000110110001;
		correct = 32'b11100101111100010011000110110001;
		#500; //-473.49695 * -1.4237587e+23 = -1.4237587e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101010100010010010011010010001;
		x2 = 32'b10010110101001010101001110111100;
		correct = 32'b01101010100010010010011010010001;
		#500; //8.290248e+25 * -2.6710032e-25 = 8.290248e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101101101100010110111010101010;
		x2 = 32'b01101010100001100000101000110000;
		correct = 32'b01101101101100111000011011010011;
		#500; //6.864079e+27 * 8.102208e+25 = 6.945101e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101101100111011110011011111;
		x2 = 32'b01011100010010100001101010100000;
		correct = 32'b01110101101100111011110011011111;
		#500; //4.556894e+32 * 2.2754888e+17 = 4.556894e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110000011101000000111101010010;
		x2 = 32'b00010101001111011011101101010010;
		correct = 32'b10110000011101000000111101010010;
		#500; //-8.8788454e-10 * 3.8316016e-26 = -8.8788454e-10
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101100010110011101010100110;
		x2 = 32'b11111111011001101110111011111010;
		correct = 32'b11111111011001101110111011111010;
		#500; //-2.4152398e-16 * -3.0696328e+38 = -3.0696328e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100000101111111101111111100;
		x2 = 32'b00111101000100010001111111001011;
		correct = 32'b11111100000101111111101111111100;
		#500; //-3.1565907e+36 * 0.03543071 = -3.1565907e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101100111111111010001011011;
		x2 = 32'b00011010010001011011100101110110;
		correct = 32'b00111101100111111111010001011011;
		#500; //0.07810279 * 4.088846e-23 = 0.07810279
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011010000001011011011111011110;
		x2 = 32'b11001110110010101111001111001101;
		correct = 32'b01011010000001011011011111011100;
		#500; //9409584000000000.0 * -1702487700.0 = 9409582000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011100111101110111110010001111;
		x2 = 32'b10110000111110110101000011101110;
		correct = 32'b10110000111110110101000011101110;
		#500; //1.6377287e-21 * -1.8285655e-09 = -1.8285655e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010001111000010000010110100110;
		x2 = 32'b01110111111110000000101011010101;
		correct = 32'b01110111111110000000101011010101;
		#500; //-3.5502222e-28 * 1.00617916e+34 = 1.00617916e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011100111001000000011011101110;
		x2 = 32'b10111110010010010111101110101000;
		correct = 32'b11011100111001000000011011101110;
		#500; //-5.134713e+17 * -0.19676077 = -5.134713e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001111111101101000001011111100;
		x2 = 32'b10011100110011010001011100010011;
		correct = 32'b01001111111101101000001011111100;
		#500; //8271558700.0 * -1.3571727e-21 = 8271558700.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011001100011000111111110111100;
		x2 = 32'b00101100100011110000000010000100;
		correct = 32'b11011001100011000111111110111100;
		#500; //-4943368000000000.0 * 4.0643617e-12 = -4943368000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110001000011001111011001001010;
		x2 = 32'b01101100100100111110001001111100;
		correct = 32'b01101100100100111110001001111100;
		#500; //-2.051268e-09 * 1.4302531e+27 = 1.4302531e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110101010011010000111111111001;
		x2 = 32'b10100110001110111010011010010110;
		correct = 32'b11110101010011010000111111111001;
		#500; //-2.5994747e+32 * -6.5104424e-16 = -2.5994747e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000110001000011111110010000010;
		x2 = 32'b00011000001110100100101101000110;
		correct = 32'b11000110001000011111110010000010;
		#500; //-10367.127 * 2.407794e-24 = -10367.127
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110000000000111101111000110011;
		x2 = 32'b00101100111001010010001111111111;
		correct = 32'b01110000000000111101111000110011;
		#500; //1.6324463e+29 * 6.512568e-12 = 1.6324463e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100110111001101101100010001;
		x2 = 32'b00010010001011111101111001001110;
		correct = 32'b10111100110111001101101100010001;
		#500; //-0.026959928 * 5.5494275e-28 = -0.026959928
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001001101110010101111011100;
		x2 = 32'b10011110011101101110001001111010;
		correct = 32'b10011110011101101110001001111010;
		#500; //-3.364326e-38 * -1.3069966e-20 = -1.3069966e-20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011011101110000011111111001101;
		x2 = 32'b01110001000100111101001011010000;
		correct = 32'b01110001000100111101001011010000;
		#500; //3.0481477e-22 * 7.3198645e+29 = 7.3198645e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011010011100000010010110100000;
		x2 = 32'b00110111001100010011000010100100;
		correct = 32'b11011010011100000010010110100000;
		#500; //-1.6898841e+16 * 1.0561347e-05 = -1.6898841e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101011101011000100011011110101;
		x2 = 32'b01100001011010100100001010011111;
		correct = 32'b01100001011010100100001010011111;
		#500; //1.224103e-12 * 2.7008367e+20 = 2.7008367e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001001001001001100001001111100;
		x2 = 32'b10101101111000110110011000111111;
		correct = 32'b01001001001001001100001001111100;
		#500; //674855.75 * -2.5852319e-11 = 674855.75
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010101001011111100110111100110;
		x2 = 32'b11000011011001100100110011001000;
		correct = 32'b11010101001011111100110111100110;
		#500; //-12081179000000.0 * -230.29993 = -12081179000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100010110000110101111101111000;
		x2 = 32'b01101000010000101111101110110100;
		correct = 32'b01101000010000101111101110110100;
		#500; //-5.2955937e-18 * 3.6831288e+24 = 3.6831288e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110010000111001000110000100010;
		x2 = 32'b00010111111101100001011011001011;
		correct = 32'b01110010000111001000110000100010;
		#500; //3.1007406e+30 * 1.5903131e-24 = 3.1007406e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111111111010000000110001110111;
		x2 = 32'b01111011111000001101010011111001;
		correct = 32'b01111011111000001101010011111001;
		#500; //1.8128804 * 2.3347882e+36 = 2.3347882e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000100100000100111010011011001;
		x2 = 32'b01110001011111101010110000100100;
		correct = 32'b01110001011111101010110000100100;
		#500; //-1043.6515 * 1.2610768e+30 = 1.2610768e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010110010101000110000111000000;
		x2 = 32'b11001100111101101110011000001100;
		correct = 32'b11010110010101000110000111011111;
		#500; //-58379075000000.0 * -129445980.0 = -58379205000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111110110101111001001011100000;
		x2 = 32'b10011110101011111111100111000100;
		correct = 32'b10111110110101111001001011100000;
		#500; //-0.42104244 * -1.8632146e-20 = -0.42104244
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110001011011101101000111101100;
		x2 = 32'b11000110111000010010001000001110;
		correct = 32'b11000110111000010010001000001110;
		#500; //-3.4752885e-09 * -28817.027 = -28817.027
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101100100010010110001001000;
		x2 = 32'b00000011110001011001011001100000;
		correct = 32'b00110101100100010010110001001000;
		#500; //1.0816229e-06 * 1.1613144e-36 = 1.0816229e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011011101010010010101001110;
		x2 = 32'b01000000000101010000001000001101;
		correct = 32'b01001011011101010010010101010000;
		#500; //16065870.0 * 2.3282502 = 16065872.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011110011001011000000001000111;
		x2 = 32'b00000001000100010001110111110101;
		correct = 32'b11011110011001011000000001000111;
		#500; //-4.134324e+18 * 2.6653787e-38 = -4.134324e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001111001101001001100111111111;
		x2 = 32'b01011011000110111101111010110111;
		correct = 32'b01011011000110111101111010110111;
		#500; //-8.904344e-30 * 4.38735e+16 = 4.38735e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100101100011011011111000100110;
		x2 = 32'b00011110101010010100100000110110;
		correct = 32'b00100101100011011100000011001011;
		#500; //2.458845e-16 * 1.7923437e-20 = 2.4590243e-16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011010001010000001110101111100;
		x2 = 32'b11001010001111111011100001011111;
		correct = 32'b11011010001010000001110101111100;
		#500; //-1.1830054e+16 * -3141143.8 = -1.1830054e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111111001010101101110110000;
		x2 = 32'b00100111101111010000000111110111;
		correct = 32'b10111111111001010101101110110000;
		#500; //-1.7918606 * 5.246017e-15 = -1.7918606
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001001100111110000110110101111;
		x2 = 32'b00110011110101010111000111010001;
		correct = 32'b11001001100111110000110110101111;
		#500; //-1302965.9 * 9.9392885e-08 = -1302965.9
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100000000001101101001100011;
		x2 = 32'b01001110110110111010101011111000;
		correct = 32'b01001110110110111010101011111000;
		#500; //-4.2633906e-22 * 1842707500.0 = 1842707500.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101001011101111100000000011;
		x2 = 32'b01101100011111010001011111110000;
		correct = 32'b01101100011111010001011111110000;
		#500; //8.226993e-36 * 1.2238851e+27 = 1.2238851e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010100101111001100001111110111;
		x2 = 32'b01111101101001011010010001001011;
		correct = 32'b01111101101001011010010001001011;
		#500; //1.9060443e-26 * 2.752196e+37 = 2.752196e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101101110011000011011111101100;
		x2 = 32'b10101000001000010010000111101000;
		correct = 32'b10101101110011000100110000010000;
		#500; //-2.321695e-11 * -8.944648e-15 = -2.3225893e-11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001101010111001111001001110;
		x2 = 32'b10110101010101111001100011101010;
		correct = 32'b10110101010101111001100011101001;
		#500; //7.621387e-14 * -8.031626e-07 = -8.0316255e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100111110101000011101011110000;
		x2 = 32'b01111001100111111110011000101010;
		correct = 32'b01111001100111111110011000101010;
		#500; //-2.0044578e+24 * 1.0378044e+35 = 1.0378044e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000010000110111010000000000010;
		x2 = 32'b01110110000100000100100111010100;
		correct = 32'b01110110000100000100100111010100;
		#500; //-1.1433522e-37 * 7.316291e+32 = 7.316291e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000010110101101010111001111101;
		x2 = 32'b01110011110100111111100000000010;
		correct = 32'b01110011110100111111100000000010;
		#500; //3.1544625e-37 * 3.3587794e+31 = 3.3587794e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000111011010011100001110011;
		x2 = 32'b10110000111111010001000001110000;
		correct = 32'b10110000111111010001000001110000;
		#500; //-6.1320063e-24 * -1.8412845e-09 = -1.8412845e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110101110111100100010000100111;
		x2 = 32'b11101000100001010101011000110000;
		correct = 32'b11101000100001010101011000110000;
		#500; //-1.6560124e-06 * -5.037317e+24 = -5.037317e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100010001101110000010000110;
		x2 = 32'b01001110011110000100101011100001;
		correct = 32'b01001110011110000100101011100001;
		#500; //-6.5802894e-22 * 1041414200.0 = 1041414200.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110110011110100001110111111010;
		x2 = 32'b10010111101001011110101111010010;
		correct = 32'b00110110011110100001110111111010;
		#500; //3.7270352e-06 * -1.07224045e-24 = 3.7270352e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011101100111001010000101010100;
		x2 = 32'b01000110111100110100000000010111;
		correct = 32'b01011101100111001010000101010100;
		#500; //1.4107993e+18 * 31136.045 = 1.4107993e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011010010100101110010001100000;
		x2 = 32'b11001010011010000001111100100100;
		correct = 32'b11001010011010000001111100100100;
		#500; //4.3611462e-23 * -3803081.0 = -3803081.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111000110101111111010100001001;
		x2 = 32'b00110011101100010001000100100011;
		correct = 32'b01111000110101111111010100001001;
		#500; //3.5041054e+34 * 8.245322e-08 = 3.5041054e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110011011110000110111111111101;
		x2 = 32'b11010100011111000111001110000101;
		correct = 32'b11010100011111000111001110000101;
		#500; //5.7843852e-08 * -4337079400000.0 = -4337079400000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000011011101110101001000100100;
		x2 = 32'b10110001100100111110010101000010;
		correct = 32'b10110001100100111110010101000010;
		#500; //7.268107e-37 * -4.3043267e-09 = -4.3043267e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101101111110001100100111001011;
		x2 = 32'b00110001000100111101101110001101;
		correct = 32'b11101101111110001100100111001011;
		#500; //-9.6245294e+27 * 2.1516116e-09 = -9.6245294e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000101001010101110010110011110;
		x2 = 32'b11000001000011011111001111000001;
		correct = 32'b11000001000011011111001111000001;
		#500; //-8.0355356e-36 * -8.87201 = -8.87201
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011110111010100011011010110000;
		x2 = 32'b11101101111111011011001110110111;
		correct = 32'b11101101111111011011001110110111;
		#500; //8.438435e+18 * -9.814621e+27 = -9.814621e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010110100101111000001110011001;
		x2 = 32'b01100001000001000010101011010110;
		correct = 32'b01100001000001000010101011010110;
		#500; //-2.4478416e-25 * 1.5237855e+20 = 1.5237855e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100101010100101101000101001;
		x2 = 32'b01101101000011101001111101011000;
		correct = 32'b01101101000011101001111101011000;
		#500; //-5853256600000.0 * 2.758719e+27 = 2.758719e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001100100000111111100000101;
		x2 = 32'b11011110000101111011110001000100;
		correct = 32'b11100001100100011010111001111110;
		#500; //-3.331855e+20 * -2.7334222e+18 = -3.3591892e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100101000011011011011110111;
		x2 = 32'b11011010000111011110011101011011;
		correct = 32'b11011010000111011110011101011011;
		#500; //-4.5962084e-12 * -1.1111487e+16 = -1.1111487e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011011101001111011111111111000;
		x2 = 32'b01111110000010010000101100000001;
		correct = 32'b01111110000010010000101100000001;
		#500; //-2.775189e-22 * 4.5540343e+37 = 4.5540343e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000100011100110001000101111110;
		x2 = 32'b11110101111000101001100011110010;
		correct = 32'b11110101111000101001100011110010;
		#500; //2.8572545e-36 * -5.7449277e+32 = -5.7449277e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100101111000111010110011100000;
		x2 = 32'b11110001010011011110011000110001;
		correct = 32'b11110001010011011110011000101111;
		#500; //1.3439577e+23 * -1.0195634e+30 = -1.0195632e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010001100011011001000110101011;
		x2 = 32'b01011101100111000001100100100010;
		correct = 32'b01011101100111000001100100100010;
		#500; //2.2335652e-28 * 1.4060074e+18 = 1.4060074e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001110101100100011001010100010;
		x2 = 32'b00011100100001101011111100100100;
		correct = 32'b11001110101100100011001010100010;
		#500; //-1494831400.0 * 8.916785e-22 = -1494831400.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001011001011101111101001010000;
		x2 = 32'b11000110000000010000111010000011;
		correct = 32'b11001011001011110001101010010100;
		#500; //-11467344.0 * -8259.628 = -11475604.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110110001010010110000011010111;
		x2 = 32'b01011001011110001110110110100101;
		correct = 32'b01011001011110001110110110100101;
		#500; //2.523933e-06 * 4379193000000000.0 = 4379193000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110000000110011011111000011100;
		x2 = 32'b11101001011000101111101110000010;
		correct = 32'b01110000000110011011101010010000;
		#500; //1.9032414e+29 * -1.7150309e+25 = 1.9030699e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101010010000011101011110011110;
		x2 = 32'b10101011000001111000101101110010;
		correct = 32'b11101010010000011101011110011110;
		#500; //-5.8585227e+25 * -4.8155154e-13 = -5.8585227e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000110010101000100111110110100;
		x2 = 32'b11111100000001110000111100101111;
		correct = 32'b11111100000001110000111100101111;
		#500; //-13587.926 * -2.805072e+36 = -2.805072e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100100101001000000110001101111;
		x2 = 32'b00100100011111101010010010011010;
		correct = 32'b01100100101001000000110001101111;
		#500; //2.4209296e+22 * 5.5216893e-17 = 2.4209296e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011001111000111110101111001000;
		x2 = 32'b00000100110000101101101100111011;
		correct = 32'b11011001111000111110101111001000;
		#500; //-8019258000000000.0 * 4.5810512e-36 = -8019258000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000110101010100100101100001100;
		x2 = 32'b01001001101100010001100011000010;
		correct = 32'b01001001101100111100000111101110;
		#500; //21797.523 * 1450776.2 = 1472573.8
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001100001101100110110111100;
		x2 = 32'b01111111010000101010010000111011;
		correct = 32'b01111111010000101010010000111011;
		#500; //-4.951904e-38 * 2.5872296e+38 = 2.5872296e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110010110110111000110010001001;
		x2 = 32'b10100010011111100100000110110100;
		correct = 32'b00110010110110111000110010001001;
		#500; //2.5558863e-08 * -3.4458202e-18 = 2.5558863e-08
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000001101001111011110111011;
		x2 = 32'b10001101001100101101110011011101;
		correct = 32'b01010000001101001111011110111011;
		#500; //12144537000.0 * -5.511634e-31 = 12144537000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100000111001110111100111111101;
		x2 = 32'b10001100001000011111011010001101;
		correct = 32'b10100000111001110111100111111101;
		#500; //-3.9213647e-19 * -1.2477183e-31 = -3.9213647e-19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110110111010101010001110100;
		x2 = 32'b00110110011001111110100001111010;
		correct = 32'b00111110110111010101010011101000;
		#500; //0.43228495 * 3.4557002e-06 = 0.4322884
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000111000110001000000101010110;
		x2 = 32'b01001001100011000000001101001111;
		correct = 32'b01001001100100001100011101011010;
		#500; //39041.336 * 1146985.9 = 1186027.2
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000110101001000100001110010100;
		x2 = 32'b10111100100111010101011011101011;
		correct = 32'b10111100100111010101011011101011;
		#500; //-6.178924e-35 * -0.019206485 = -0.019206485
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010110101000001000100111110001;
		x2 = 32'b01110101110000000000100110001001;
		correct = 32'b01110101110000000000100110001001;
		#500; //2.5936447e-25 * 4.8687226e+32 = 4.8687226e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001111100110100001101001000;
		x2 = 32'b11000010000011100000100001001011;
		correct = 32'b11000010100000111101010011111000;
		#500; //-30.407852 * -35.5081 = -65.915955
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111001000110111111001101110110;
		x2 = 32'b00011100010111110011101100000110;
		correct = 32'b10111001000110111111001101110110;
		#500; //-0.00014872648 * 7.3860797e-22 = -0.00014872648
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010010111011001000100110010111;
		x2 = 32'b01101001100111100111000011111000;
		correct = 32'b01101001100111100111000011111000;
		#500; //507960330000.0 * 2.394297e+25 = 2.394297e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110110111001000101111110010000;
		x2 = 32'b10110100100111010100111011110100;
		correct = 32'b11110110111001000101111110010000;
		#500; //-2.3159803e+33 * -2.9300975e-07 = -2.3159803e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100001000010101000000110101110;
		x2 = 32'b01010011000010101000111010101101;
		correct = 32'b01010011000010101000111010101101;
		#500; //-4.692785e-19 * 595099200000.0 = 595099200000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110001001111000010011010010100;
		x2 = 32'b11011001100011011001100110011010;
		correct = 32'b01110001001111000010011010010100;
		#500; //9.316771e+29 * -4982107300000000.0 = 9.316771e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101110010111100000001000000001;
		x2 = 32'b01000101011000000011111011000000;
		correct = 32'b01000101011000000011111011000000;
		#500; //5.0478736e-11 * 3587.9219 = 3587.9219
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000101100001101101111100111111;
		x2 = 32'b00010001011000101110110100001011;
		correct = 32'b01000101100001101101111100111111;
		#500; //4315.906 * 1.7901301e-28 = 4315.906
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110001101001000101111111001011;
		x2 = 32'b11101110011010010101001111001011;
		correct = 32'b11101110011010010101001111001011;
		#500; //4.7839186e-09 * -1.8052827e+28 = -1.8052827e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001001111010100010111001111001;
		x2 = 32'b10011000001100110011011100010000;
		correct = 32'b01001001111010100010111001111001;
		#500; //1918415.1 * -2.3163007e-24 = 1918415.1
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110010010011011000000000000000;
		x2 = 32'b11001101110101110001001001111001;
		correct = 32'b01110010010011011000000000000000;
		#500; //4.070347e+30 * -451039000.0 = 4.070347e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100100000111101101000000100;
		x2 = 32'b10001010100100011000011101000111;
		correct = 32'b10010100100000111101101000001101;
		#500; //-1.3313612e-26 * -1.4013878e-32 = -1.3313626e-26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010110101111010110100110110011;
		x2 = 32'b10010000000011111010000001110110;
		correct = 32'b00010110101111010110010100110110;
		#500; //3.0601302e-25 * -2.8325392e-29 = 3.059847e-25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110011011111001111111001110001;
		x2 = 32'b11111001100111100000110111000100;
		correct = 32'b11111001100111100001010110101100;
		#500; //-2.0044243e+31 * -1.0258276e+35 = -1.0260281e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111110000100100000110001101;
		x2 = 32'b10010110001100110101010011100011;
		correct = 32'b11111111110000100100000110001101;
		#500; //nan * -1.448629e-25 = nan
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100111001100110111110000110001;
		x2 = 32'b10101001100001011000101110111100;
		correct = 32'b11100111001100110111110000110001;
		#500; //-8.475945e+23 * -5.9306265e-14 = -8.475945e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001010011100000100111110101001;
		x2 = 32'b00010111001000010110101100111110;
		correct = 32'b11001010011100000100111110101001;
		#500; //-3937258.2 * 5.2157264e-25 = -3937258.2
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011101010010000101111000001101;
		x2 = 32'b10110000000010010101000011001011;
		correct = 32'b11011101010010000101111000001101;
		#500; //-9.023745e+17 * -4.9955123e-10 = -9.023745e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011001001110101011110110001110;
		x2 = 32'b00111011100110110101100011111001;
		correct = 32'b00111011100110110101100011111001;
		#500; //-9.654255e-24 * 0.004740831 = 0.004740831
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001100011100001000001101001011;
		x2 = 32'b01111010110101100001011111100101;
		correct = 32'b01111010110101100001011111100101;
		#500; //-63049004.0 * 5.558181e+35 = 5.558181e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101101000111111000111101000;
		x2 = 32'b00010011100100001110110010000000;
		correct = 32'b01111101101000111111000111101000;
		#500; //2.7240027e+37 * 3.6583918e-27 = 2.7240027e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011000110001001100111100111001;
		x2 = 32'b00000000100110111110110100010101;
		correct = 32'b00011000110001001100111100111001;
		#500; //5.0874054e-24 * 1.4319551e-38 = 5.0874054e-24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101010001111110111110110011111;
		x2 = 32'b01110110011010110001011010110001;
		correct = 32'b01110110011010110001011010110000;
		#500; //-5.7874515e+25 * 1.192041e+33 = 1.1920409e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110000011100100100011111110011;
		x2 = 32'b10001111101011101000100101100101;
		correct = 32'b01110000011100100100011111110011;
		#500; //2.9992941e+29 * -1.7210647e-29 = 2.9992941e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001011100100000111111111010;
		x2 = 32'b11011010010100001010100110110111;
		correct = 32'b11011010010100001010100110110111;
		#500; //-15.128901 * -1.468335e+16 = -1.468335e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100001110111000001001010010111;
		x2 = 32'b00010010110101010101101110010101;
		correct = 32'b01100001110111000001001010010111;
		#500; //5.074529e+20 * 1.3464767e-27 = 5.074529e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010100110010001001110000101;
		x2 = 32'b00001001001101000000110000111110;
		correct = 32'b01000010100110010001001110000101;
		#500; //76.538124 * 2.1672468e-33 = 76.538124
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001001010011101110001110010001;
		x2 = 32'b10010001011110111110011000100010;
		correct = 32'b10010001011110111110011011110001;
		#500; //-2.490335e-33 * -1.9871324e-28 = -1.9871573e-28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011000011010101101100001101;
		x2 = 32'b01111101101011011001101010100011;
		correct = 32'b01111101101011011001101010100011;
		#500; //-4.1540697e-37 * 2.884492e+37 = 2.884492e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100111000011000101101110001011;
		x2 = 32'b11010110010100100100010110111011;
		correct = 32'b11100111000011000101101110001011;
		#500; //-6.6282e+23 * -57799233000000.0 = -6.6282e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110001000101101100111000001010;
		x2 = 32'b01101010001010100111010101110010;
		correct = 32'b01110001000101101101000010110100;
		#500; //7.467494e+29 * 5.1518e+25 = 7.468009e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101100001000100110110010101001;
		x2 = 32'b11110010111100010010100100010011;
		correct = 32'b11110010111100010010100100010011;
		#500; //2.3081903e-12 * -9.5533495e+30 = -9.5533495e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110101010110110100101111100010;
		x2 = 32'b11011110011001001111100010101100;
		correct = 32'b11011110011001001111100010101100;
		#500; //-8.169428e-07 * -4.1247816e+18 = -4.1247816e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000000100010010001101011001011;
		x2 = 32'b00000111111000100010110000011001;
		correct = 32'b00000111111000100010100111110101;
		#500; //-1.2591074e-38 * 3.403062e-34 = 3.402936e-34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111111110010010000000000000;
		x2 = 32'b10011101001000001110000101110110;
		correct = 32'b10111111111110010010000000000000;
		#500; //-1.9462891 * -2.1292384e-21 = -1.9462891
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000110111010011101101001111000;
		x2 = 32'b10000011101101011111000101110101;
		correct = 32'b10000110111011001011001000111110;
		#500; //-8.796587e-35 * -1.069366e-36 = -8.9035237e-35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101100000001101000110010010110;
		x2 = 32'b10000000001110111001100100111111;
		correct = 32'b00101100000001101000110010010110;
		#500; //1.9120586e-12 * -5.473269e-39 = 1.9120586e-12
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001100100100010010000010000;
		x2 = 32'b10110111111010111010111110010100;
		correct = 32'b11000001100100100010010000011111;
		#500; //-18.267609 * -2.8095943e-05 = -18.267637
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011100110100101010010101111;
		x2 = 32'b00011100001000000100010010010101;
		correct = 32'b01101011100110100101010010101111;
		#500; //3.7314897e+26 * 5.30282e-22 = 3.7314897e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110001010000010110000000011;
		x2 = 32'b01101110011100101100111000110001;
		correct = 32'b01101110011100101100111000110001;
		#500; //-3.8237868e-11 * 1.8786161e+28 = 1.8786161e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000000100001110010100000111111;
		x2 = 32'b10011110111101010001111111011101;
		correct = 32'b11000000100001110010100000111111;
		#500; //-4.223663 * -2.5953562e-20 = -4.223663
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001010000110100001000100101111;
		x2 = 32'b00101001001000010100001001010001;
		correct = 32'b01001010000110100001000100101111;
		#500; //2524235.8 * 3.5806702e-14 = 2524235.8
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101000000000100111110101010001;
		x2 = 32'b01000001011101010110011101011101;
		correct = 32'b11101000000000100111110101010001;
		#500; //-2.4648773e+24 * 15.337735 = -2.4648773e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101011110010011110111101101011;
		x2 = 32'b10110001100101100010011010001001;
		correct = 32'b10110001100101100011001100101000;
		#500; //-1.4348361e-12 * -4.3699555e-09 = -4.3713904e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110000010001001001010111001101;
		x2 = 32'b01011000110001011100110001001111;
		correct = 32'b01011000110001011100110001001111;
		#500; //-7.1517264e-10 * 1739850300000000.0 = 1739850300000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111001001101111001100011100010;
		x2 = 32'b00101101101001010100001011100101;
		correct = 32'b11111001001101111001100011100010;
		#500; //-5.9580697e+34 * 1.8788035e-11 = -5.9580697e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101001111000010010100010010011;
		x2 = 32'b11001100100011010010101001100000;
		correct = 32'b01101001111000010010100010010011;
		#500; //3.402499e+25 * -74011390.0 = 3.402499e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001100011110111111001010111101;
		x2 = 32'b00011100110000011011011100000000;
		correct = 32'b00011100110000011011011100000000;
		#500; //-1.9409383e-31 * 1.2818973e-21 = 1.2818973e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110011100111100001110010111111;
		x2 = 32'b00011000111110001100111010000011;
		correct = 32'b01110011100111100001110010111111;
		#500; //2.5053892e+31 * 6.431502e-24 = 2.5053892e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101110101001000011100101001000;
		x2 = 32'b00000101100001100000100100000111;
		correct = 32'b00101110101001000011100101001000;
		#500; //7.468032e-11 * 1.2604616e-35 = 7.468032e-11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100001110000011000100001010111;
		x2 = 32'b10111101000001001100111001010011;
		correct = 32'b10111101000001001100111001010011;
		#500; //-1.3114278e-18 * -0.03242333 = -0.03242333
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100010100001111001101000000101;
		x2 = 32'b01000111100001100110111110001000;
		correct = 32'b01100010100001111001101000000101;
		#500; //1.2507044e+21 * 68831.06 = 1.2507044e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110110111100010111010100101101;
		x2 = 32'b01111110111100010010101010111101;
		correct = 32'b01111110111100010010101010111101;
		#500; //7.1960008e-06 * 1.6028293e+38 = 1.6028293e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110100110000010001100110000100;
		x2 = 32'b00010000101011100010011000111001;
		correct = 32'b10110100110000010001100110000100;
		#500; //-3.5967616e-07 * 6.868979e-29 = -3.5967616e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110100111101010111010000011000;
		x2 = 32'b10000101001001111100001111101001;
		correct = 32'b10110100111101010111010000011000;
		#500; //-4.5719275e-07 * -7.888285e-36 = -4.5719275e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111001010001011100011100000011;
		x2 = 32'b11010110100010111101001010000110;
		correct = 32'b11111001010001011100011100000011;
		#500; //-6.418243e+34 * -76868150000000.0 = -6.418243e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010110100110000010001110010001;
		x2 = 32'b10100111111001101100111101010001;
		correct = 32'b10100111111001101100111101010001;
		#500; //2.457937e-25 * -6.4062597e-15 = -6.4062597e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101110101000110101110111101111;
		x2 = 32'b01110000000110110101101010010011;
		correct = 32'b01110000000001101110111011010101;
		#500; //-2.5279808e+28 * 1.923187e+29 = 1.6703889e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010110000100000100110111010100;
		x2 = 32'b10001111001100000001010100101111;
		correct = 32'b01010110000100000100110111010100;
		#500; //39665986000000.0 * -8.68155e-30 = 39665986000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001101001110101101111111000011;
		x2 = 32'b10111011011110110011001001111001;
		correct = 32'b10111011011110110011001001111001;
		#500; //-5.758502e-31 * -0.0038329645 = -0.0038329645
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110101100000000101000110011000;
		x2 = 32'b01101100001011100111000110000001;
		correct = 32'b11110101100000000101000110000010;
		#500; //-3.253266e+32 * 8.435564e+26 = -3.2532577e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010010000011100000110011100011;
		x2 = 32'b11100110110100101011000001110111;
		correct = 32'b11100110110100101011000001110111;
		#500; //-152525390000.0 * -4.9747608e+23 = -4.9747608e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100111100001010100010110001101;
		x2 = 32'b11001001011110001110010001001001;
		correct = 32'b11001001011110001110010001001001;
		#500; //-3.6990323e-15 * -1019460.56 = -1019460.56
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111001010110011000110001111;
		x2 = 32'b01000100111001000000101111110010;
		correct = 32'b01000100111001000000101111110010;
		#500; //2.3757883e-15 * 1824.3733 = 1824.3733
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111100110111010110111111011;
		x2 = 32'b00110011101010101110110000010111;
		correct = 32'b10110111100110110000001100001111;
		#500; //-1.8558456e-05 * 7.9591864e-08 = -1.8478864e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011011011001100011111011111;
		x2 = 32'b11100111110101111111100110111101;
		correct = 32'b11100111110101111111100110111101;
		#500; //-6.9583607e-37 * -2.0398313e+24 = -2.0398313e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100101111010010110010101101000;
		x2 = 32'b11000111000111111001000111010000;
		correct = 32'b11000111000111111001000111010000;
		#500; //4.0487773e-16 * -40849.812 = -40849.812
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100000110110011011010000010;
		x2 = 32'b01101001001010011110000100000100;
		correct = 32'b01101001001010011110000100000100;
		#500; //-7.83625e-27 * 1.2835692e+25 = 1.2835692e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110000001100100100101011001111;
		x2 = 32'b11010110100111010100110111011100;
		correct = 32'b11010110100111010100110111011100;
		#500; //6.486233e-10 * -86478865000000.0 = -86478865000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110010100110011110000111011110;
		x2 = 32'b10000000000000000001000100101001;
		correct = 32'b11110010100110011110000111011110;
		#500; //-6.0959057e+30 * -6.156e-42 = -6.0959057e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110011100010001000010111000110;
		x2 = 32'b10100110000000111101011000000011;
		correct = 32'b11110011100010001000010111000110;
		#500; //-2.1632862e+31 * -4.5739795e-16 = -2.1632862e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100111111010101101101001000;
		x2 = 32'b10110001001000010010010100110101;
		correct = 32'b00111100111111010101101101000111;
		#500; //0.030927315 * -2.3449733e-09 = 0.030927313
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010001000000101010101011101101;
		x2 = 32'b11001011110011010111011001011100;
		correct = 32'b11001011110011010111011001011100;
		#500; //1.0307862e-28 * -26930360.0 = -26930360.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010001101001111000110011001000;
		x2 = 32'b11110010111110100100000101001100;
		correct = 32'b11110010111110100100000101001100;
		#500; //2.6434717e-28 * -9.9136245e+30 = -9.9136245e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111110010110100110110111000;
		x2 = 32'b01000101000111011111110110110110;
		correct = 32'b11011111110010110100110110111000;
		#500; //-2.9299135e+19 * 2527.857 = -2.9299135e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001110001100010101000100110001;
		x2 = 32'b00100010111100110001001010000011;
		correct = 32'b11001110001100010101000100110001;
		#500; //-743722050.0 * 6.588488e-18 = -743722050.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011101000110010100110101000001;
		x2 = 32'b10001011101100011000111111010010;
		correct = 32'b10011101000110010100110101000001;
		#500; //-2.028932e-21 * -6.8394317e-32 = -2.028932e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000000100111001101110000001110;
		x2 = 32'b00011010111010101100010110100010;
		correct = 32'b00011010111010101100010110100010;
		#500; //-1.4405278e-38 * 9.7099425e-23 = 9.7099425e-23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001110011100000101100010100001;
		x2 = 32'b00011010101111101110001010000010;
		correct = 32'b01001110011100000101100010100001;
		#500; //1008085060.0 * 7.89481e-23 = 1008085060.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101011100100110100010011111010;
		x2 = 32'b10110101101100000010100001001101;
		correct = 32'b10110101101100000010100001000100;
		#500; //1.0464123e-12 * -1.3124751e-06 = -1.3124741e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010010010010010110100001001;
		x2 = 32'b10010001110101101111111100101100;
		correct = 32'b01000010010010010010110100001001;
		#500; //50.29398 * -3.3920509e-28 = 50.29398
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100111010000100111101001000;
		x2 = 32'b10000101110001110010101011101110;
		correct = 32'b01110100111010000100111101001000;
		#500; //1.4724376e+32 * -1.872964e-35 = 1.4724376e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100100001000011011110001010111;
		x2 = 32'b00001000000011001111001100101111;
		correct = 32'b11100100001000011011110001010111;
		#500; //-1.1933988e+22 * 4.241558e-34 = -1.1933988e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110010101110101011101000011;
		x2 = 32'b01100010001000100011001111110010;
		correct = 32'b01100010001000100011001111110010;
		#500; //-3.208829e-06 * 7.480289e+20 = 7.480289e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110001111010010101000101010011;
		x2 = 32'b10000111111110001011110000101010;
		correct = 32'b11110001111010010101000101010011;
		#500; //-2.3106663e+30 * -3.7425486e-34 = -2.3106663e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001000110110010011000100000;
		x2 = 32'b11101001011110101110010100001010;
		correct = 32'b11101001011110101110010110100101;
		#500; //-1.7887453e+20 * -1.8957066e+25 = -1.8957245e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100001000000111001011101010001;
		x2 = 32'b10110100001000101111010001011111;
		correct = 32'b10110100001000101111010001011111;
		#500; //4.458479e-19 * -1.5176327e-07 = -1.5176327e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110001011010000001101000111011;
		x2 = 32'b10000011000111100111000000101010;
		correct = 32'b10110001011010000001101000111011;
		#500; //-3.3775354e-09 * -4.6560785e-37 = -3.3775354e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011111000110011100100101101;
		x2 = 32'b00111000111100000111111001100110;
		correct = 32'b01001011111000110011100100101101;
		#500; //29782618.0 * 0.00011467635 = 29782618.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110010111101001001101110110;
		x2 = 32'b11001011010010011110001110110101;
		correct = 32'b11001011010010011110001110110101;
		#500; //-5.0607928e-11 * -13231029.0 = -13231029.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010101001111100000111111111001;
		x2 = 32'b10010010100111110001101100110010;
		correct = 32'b11010101001111100000111111111001;
		#500; //-13060988000000.0 * -1.0041015e-27 = -13060988000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011101110101010101011100101;
		x2 = 32'b10110010100101000011000111011010;
		correct = 32'b11111011101110101010101011100101;
		#500; //-1.9384667e+36 * -1.7252137e-08 = -1.9384667e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000110011011011111011010011;
		x2 = 32'b11110110010110111000101010011001;
		correct = 32'b11110110010110111010010001010001;
		#500; //-5.0940095e+29 * -1.1132071e+33 = -1.11371655e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111001100011101011001101111111;
		x2 = 32'b10000001111011100100100001011100;
		correct = 32'b00111001100011101011001101111111;
		#500; //0.00027218086 * -8.7531223e-38 = 0.00027218086
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111111010100111100101011110011;
		x2 = 32'b11010010001101101110100000110100;
		correct = 32'b11010010001101101110100000110100;
		#500; //0.8273155 * -196394940000.0 = -196394940000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100101101100011101000101011001;
		x2 = 32'b00111101011010000101101100011111;
		correct = 32'b11100101101100011101000101011001;
		#500; //-1.0496508e+23 * 0.056727525 = -1.0496508e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011110111100100111111100000001;
		x2 = 32'b10110111010000110000110001000111;
		correct = 32'b10110111010000110000110001000111;
		#500; //2.5675274e-20 * -1.1625764e-05 = -1.1625764e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111010100001000000111000000110;
		x2 = 32'b00010110100001110000010011100101;
		correct = 32'b10111010100001000000111000000110;
		#500; //-0.001007498 * 2.1813515e-25 = -0.001007498
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110111010001111110010000110;
		x2 = 32'b00101110100000110111101011000010;
		correct = 32'b00111110111010001111110010000110;
		#500; //0.4550516 * 5.9789965e-11 = 0.4550516
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000110011000011011010001110110;
		x2 = 32'b01000110101110011010110010111100;
		correct = 32'b01000111000101010100001101111100;
		#500; //14445.115 * 23766.367 = 38211.484
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100000101000010010010001110;
		x2 = 32'b01010011011001101101011011000010;
		correct = 32'b11111100000101000010010010001110;
		#500; //-3.0768054e+36 * 991445500000.0 = -3.0768054e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111100110011101000110010011;
		x2 = 32'b10000000101010101100001011110111;
		correct = 32'b11010111100110011101000110010011;
		#500; //-338250800000000.0 * -1.5681975e-38 = -338250800000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111001101001001011011010111100;
		x2 = 32'b01111100011001110000100000011101;
		correct = 32'b01111100011001110000100000011101;
		#500; //0.00031416665 * 4.7983405e+36 = 4.7983405e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010101111011101011000000010001;
		x2 = 32'b11100011101011011100001111010110;
		correct = 32'b11100011101011011100001111010110;
		#500; //-9.640522e-26 * -6.4107964e+21 = -6.4107964e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100001100111001001001000101111;
		x2 = 32'b10011011100101100101111011000110;
		correct = 32'b01100001100111001001001000101111;
		#500; //3.610282e+20 * -2.4876664e-22 = 3.610282e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010011101111001111111001000010;
		x2 = 32'b11110100000010111000000111110011;
		correct = 32'b11110100000010111000000111110011;
		#500; //-4.770859e-27 * -4.421173e+31 = -4.421173e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100110100010000001110011111;
		x2 = 32'b10111010101010110011110010001000;
		correct = 32'b01110100110100010000001110011111;
		#500; //1.3247845e+32 * -0.0013064304 = 1.3247845e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000011100010000000001000010101;
		x2 = 32'b01100101111101011000001010000100;
		correct = 32'b01100101111101011000001010000100;
		#500; //7.99384e-37 * 1.4492342e+23 = 1.4492342e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100100001001110010000000011;
		x2 = 32'b00000100011000011001100011100101;
		correct = 32'b10101100100001001110010000000011;
		#500; //-3.77698e-12 * 2.6518829e-36 = -3.77698e-12
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101011100101001010110010100100;
		x2 = 32'b10101001001011111111101100111100;
		correct = 32'b11101011100101001010110010100100;
		#500; //-3.594726e+26 * -3.9075717e-14 = -3.594726e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110111001010001111010110000100;
		x2 = 32'b11001101110110010100010100100001;
		correct = 32'b11110111001010001111010110000100;
		#500; //-3.4268966e+33 * -455648300.0 = -3.4268966e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100111101001000010110100111010;
		x2 = 32'b01100101101001000011110110011011;
		correct = 32'b01100101101001000011110110011011;
		#500; //-4.556818e-15 * 9.6950565e+22 = 9.6950565e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000101001010010011001010001100;
		x2 = 32'b10111110011110010011011101000000;
		correct = 32'b10111110011110010011011101000000;
		#500; //-7.955626e-36 * -0.24337482 = -0.24337482
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110010101001101100000110100;
		x2 = 32'b00010100100100111010110010111011;
		correct = 32'b00111110010101001101100000110100;
		#500; //0.207856 * 1.4911337e-26 = 0.207856
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010110111100100011000110000111;
		x2 = 32'b00100011111011110110010100101101;
		correct = 32'b11010110111100100011000110000111;
		#500; //-133147270000000.0 * 2.5955282e-17 = -133147270000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110111110110010111001011010101;
		x2 = 32'b10011110011010010100001001010010;
		correct = 32'b01110111110110010111001011010101;
		#500; //8.8207616e+33 * -1.2348632e-20 = 8.8207616e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000000001000100010011011110111;
		x2 = 32'b01101001011110111101010000101011;
		correct = 32'b01101001011110111101010000101011;
		#500; //-3.136385e-39 * 1.9027645e+25 = 1.9027645e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011001100101101011010001011010;
		x2 = 32'b10010100000001001110001111110011;
		correct = 32'b00011001100101101010001110111110;
		#500; //1.558248e-23 * -6.709252e-27 = 1.5575771e-23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101011110101010000001111010;
		x2 = 32'b01000000111001110001000011110101;
		correct = 32'b01000000111001110001000011110101;
		#500; //1.17844184e-35 * 7.22082 = 7.22082
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010001101001001100100110100110;
		x2 = 32'b11001110011001100100000100010000;
		correct = 32'b01010001101000101111110100100100;
		#500; //88469720000.0 * -965755900.0 = 87503960000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001100000110100111000011011010;
		x2 = 32'b01001111100101000101110001100010;
		correct = 32'b01001111100101000101110001100010;
		#500; //-1.1897688e-31 * 4978164700.0 = 4978164700.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110010011001000001010111001;
		x2 = 32'b10010101011111100010101001011111;
		correct = 32'b10101110010011001000001010111001;
		#500; //-4.6500335e-11 * -5.1328316e-26 = -4.6500335e-11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110010000011001101111100010110;
		x2 = 32'b10000010001011000101001101111011;
		correct = 32'b11110010000011001101111100010110;
		#500; //-2.790246e+30 * -1.2660522e-37 = -2.790246e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101011100100111110111111000110;
		x2 = 32'b00011111111000100110110010110110;
		correct = 32'b10101011100100111110111111000101;
		#500; //-1.0511529e-12 * 9.589457e-20 = -1.0511528e-12
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101001001010100100110000110111;
		x2 = 32'b00001100111111010000000110100001;
		correct = 32'b01101001001010100100110000110111;
		#500; //1.2867331e+25 * 3.8981802e-31 = 1.2867331e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010101100101100011111011110010;
		x2 = 32'b11000101101110110111110010100110;
		correct = 32'b11000101101110110111110010100110;
		#500; //6.068383e-26 * -5999.581 = -5999.581
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000000001101001111100001100101;
		x2 = 32'b00011100011010100000100000111011;
		correct = 32'b00011100011010100000100000111011;
		#500; //4.864553e-39 * 7.7434743e-22 = 7.7434743e-22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011101001111111000010001110111;
		x2 = 32'b00000010111100101111001001011100;
		correct = 32'b10011101001111111000010001110111;
		#500; //-2.5347122e-21 * 3.5697812e-37 = -2.5347122e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101010100010001000100010101000;
		x2 = 32'b00010000100111111111000010111100;
		correct = 32'b00101010100010001000100010101000;
		#500; //2.4253277e-13 * 6.308535e-29 = 2.4253277e-13
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100001010100000000001111100;
		x2 = 32'b10111010011110011001011111010001;
		correct = 32'b11110100001010100000000001111100;
		#500; //-5.387575e+31 * -0.00095212186 = -5.387575e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110000101111110001010101111000;
		x2 = 32'b10001000010000001101010110101011;
		correct = 32'b01110000101111110001010101111000;
		#500; //4.7310073e+29 * -5.8029064e-34 = 4.7310073e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100010101001111101011010001110;
		x2 = 32'b01000010100001110100010000000100;
		correct = 32'b01000010100001110100010000000100;
		#500; //-4.549261e-18 * 67.63284 = 67.63284
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000100011000001010110111000001;
		x2 = 32'b00000110010000010100101100001001;
		correct = 32'b00000110010011110101010111100101;
		#500; //2.6410857e-36 * 3.6354393e-35 = 3.8995478e-35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001001110111011011001010001;
		x2 = 32'b11000000011110111111101101110010;
		correct = 32'b11000001011110101011010100101110;
		#500; //-11.732011 * -3.937222 = -15.669233
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110110110011001100011000110;
		x2 = 32'b11110110011011101101100011011010;
		correct = 32'b11110110011011101101100011011010;
		#500; //-9.8951555e-11 * -1.21109856e+33 = -1.21109856e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101010101100011100100111011;
		x2 = 32'b10000110010101001101001011001100;
		correct = 32'b00110101010101100011100100111011;
		#500; //7.9804494e-07 * -4.0027637e-35 = 7.9804494e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000110110001110100010111111101;
		x2 = 32'b00000111101101011000000111010101;
		correct = 32'b01000110110001110100010111111101;
		#500; //25506.994 * 2.7310162e-34 = 25506.994
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111001001100011000011111111100;
		x2 = 32'b11110100010111011111001001111100;
		correct = 32'b11110100010111011111001001111100;
		#500; //-0.00016930694 * -7.0337877e+31 = -7.0337877e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111100001101000111011101110;
		x2 = 32'b11011101011000001011000100010101;
		correct = 32'b11011111100011011001010001110111;
		#500; //-1.9391897e+19 * -1.0119216e+18 = -2.040382e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011101010110010001010001111;
		x2 = 32'b10110000100011101011100000101001;
		correct = 32'b10110000100011101011100000101001;
		#500; //1.8554493e-17 * -1.0384201e-09 = -1.0384201e-09
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010101110010000111001011011000;
		x2 = 32'b10001101111001010011010000101001;
		correct = 32'b11010101110010000111001011011000;
		#500; //-27549447000000.0 * -1.4125772e-30 = -27549447000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001011110010101100010101011111;
		x2 = 32'b11111111010010010000101001000111;
		correct = 32'b11111111010010010000101001000111;
		#500; //-26577598.0 * -2.672282e+38 = -2.672282e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110010001010000001111110010111;
		x2 = 32'b10100101111011111110100000101101;
		correct = 32'b11110010001010000001111110010111;
		#500; //-3.330027e+30 * -4.161722e-16 = -3.330027e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110100111110000111000110001101;
		x2 = 32'b00000001011111101010111100100001;
		correct = 32'b10110100111110000111000110001101;
		#500; //-4.627622e-07 * 4.677808e-38 = -4.627622e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110011010110110100111000010;
		x2 = 32'b10101011000001101001111010010101;
		correct = 32'b10110110011010110110100111000100;
		#500; //-3.5079288e-06 * -4.782644e-13 = -3.5079293e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000001101100010011101100011;
		x2 = 32'b00111000100111011000101110011000;
		correct = 32'b00111000100111011000101110011000;
		#500; //3.5923514e-29 * 7.512345e-05 = 7.512345e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000011111111101110100001111111;
		x2 = 32'b01110100001011010000011010111100;
		correct = 32'b01110100001011010000011010111100;
		#500; //1.4982157e-36 * 5.4834225e+31 = 5.4834225e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010001000000100011010011101;
		x2 = 32'b00001000101011001101110011010101;
		correct = 32'b10101010001000000100011010011101;
		#500; //-1.4235354e-13 * 1.0403791e-33 = -1.4235354e-13
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101100011101000001101101010110;
		x2 = 32'b00000110100000111000011100100000;
		correct = 32'b11101100011101000001101101010110;
		#500; //-1.18042796e+27 * 4.947527e-35 = -1.18042796e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101100011001101101000011110001;
		x2 = 32'b00110000110000111010001001000110;
		correct = 32'b11101100011001101101000011110001;
		#500; //-1.11615855e+27 * 1.4234238e-09 = -1.11615855e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011100001110110110100110110;
		x2 = 32'b00111010100011100100101001001100;
		correct = 32'b11111011100001110110110100110110;
		#500; //-1.4063503e+36 * 0.0010855882 = -1.4063503e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111011100111100110110000011001;
		x2 = 32'b00011110111101001100101000010100;
		correct = 32'b01111011100111100110110000011001;
		#500; //1.6451508e+36 * 2.5918082e-20 = 1.6451508e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011001101011110110011110000010;
		x2 = 32'b10111100110011101001111001000000;
		correct = 32'b11011001101011110110011110000010;
		#500; //-6171491000000000.0 * -0.025221944 = -6171491000000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101100000011101010100111011010;
		x2 = 32'b01000101010000100000001001000000;
		correct = 32'b11101100000011101010100111011010;
		#500; //-6.898783e+26 * 3104.1406 = -6.898783e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010001001110101011011001101010;
		x2 = 32'b01100001101101101010101101001111;
		correct = 32'b01100001101101101010101101001111;
		#500; //50120270000.0 * 4.2120644e+20 = 4.2120644e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101010100001011100111100000101;
		x2 = 32'b11010100111000111110000000001100;
		correct = 32'b01101010100001011100111100000101;
		#500; //8.088238e+25 * -7829731700000.0 = 8.088238e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011111101111011011110100111;
		x2 = 32'b01110100100110001000110100010111;
		correct = 32'b01110100100110001000110100010111;
		#500; //-1.455952e-36 * 9.669077e+31 = 9.669077e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100010010000010001111111110;
		x2 = 32'b01000110101101110111010011111000;
		correct = 32'b11110100010010000010001111111110;
		#500; //-6.3427086e+31 * 23482.484 = -6.3427086e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010011000011000011001001000101;
		x2 = 32'b00100100100010101001101111000011;
		correct = 32'b00100100100010101001101111000011;
		#500; //1.769527e-27 * 6.011183e-17 = 6.011183e-17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100010000110100010011111010;
		x2 = 32'b11110111010011110011001110000111;
		correct = 32'b11110111010011110011001110000111;
		#500; //-6.460924e-22 * -4.2025412e+33 = -4.2025412e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010000100101100010011011011;
		x2 = 32'b10100100110100101110100101011101;
		correct = 32'b10101010000100101101111100111000;
		#500; //-1.3035703e-13 * -9.1468315e-17 = -1.304485e-13
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100010011001011110000100000101;
		x2 = 32'b00100000101100100100111011000001;
		correct = 32'b11100010011001011110000100000101;
		#500; //-1.0601297e+21 * 3.0206488e-19 = -1.0601297e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010111000011001110100001100111;
		x2 = 32'b01010001001011001010000011100010;
		correct = 32'b01010111000011001111001100110001;
		#500; //154929790000000.0 * 46339596000.0 = 154976130000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100001111000111010000100011100;
		x2 = 32'b11101000110101111000001110001011;
		correct = 32'b11101000110101110111111111111100;
		#500; //5.248775e+20 * -8.1418827e+24 = -8.1413575e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010001110111111101010111110111;
		x2 = 32'b10000011101111010100100001000001;
		correct = 32'b11010001110111111101010111110111;
		#500; //-120170930000.0 * -1.112501e-36 = -120170930000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110010111101011100111101100;
		x2 = 32'b00010100100110001000110111011110;
		correct = 32'b10110110010111101011100111101100;
		#500; //-3.3188799e-06 * 1.5404035e-26 = -3.3188799e-06
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111001011011001000101101000001;
		x2 = 32'b10110010001011101000011011011011;
		correct = 32'b00111001011011001000100010000111;
		#500; //0.0002255859 * -1.0158796e-08 = 0.00022557574
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001101001001010001111100100110;
		x2 = 32'b11110110110111011101110000100000;
		correct = 32'b11110110110111011101110000100000;
		#500; //-5.0882044e-31 * -2.2499263e+33 = -2.2499263e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111010101011101010100010000;
		x2 = 32'b11100100011000001110101110011000;
		correct = 32'b11100100011000001110101110011000;
		#500; //2.967519e-15 * -1.6596188e+22 = -1.6596188e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010000011001001110111000011;
		x2 = 32'b11111001010010001111010010110100;
		correct = 32'b11111001010010001111010010110100;
		#500; //-1.2489232e-13 * -6.521391e+34 = -6.521391e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000101000001011010111100101000;
		x2 = 32'b10001000001111111101000101010100;
		correct = 32'b11000101000001011010111100101000;
		#500; //-2138.9473 * -5.7723036e-34 = -2138.9473
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011011011010111101110010110010;
		x2 = 32'b10101011111101010011110001101110;
		correct = 32'b01011011011010111101110010110010;
		#500; //6.6389277e+16 * -1.742507e-12 = 6.6389277e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111111100011011010100110101000;
		x2 = 32'b10111100110101011100010000110100;
		correct = 32'b00111111100010100101001010010111;
		#500; //1.10674 * -0.026094534 = 1.0806454
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110010000000011110100111111;
		x2 = 32'b11001100100000000011110000011110;
		correct = 32'b11001100100000000011110000011110;
		#500; //-4.3710143e-11 * -67231980.0 = -67231980.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011101011011101110101000001011;
		x2 = 32'b10001010001111110100001111001111;
		correct = 32'b00011101011011101110101000001011;
		#500; //3.1620035e-21 * -9.209069e-33 = 3.1620035e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011001001111110011101000100001;
		x2 = 32'b11001100101011000000010101100101;
		correct = 32'b11001100101011000000010101100101;
		#500; //-9.8862076e-24 * -90188584.0 = -90188584.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101100100100100111101010011110;
		x2 = 32'b10001010100100011101100101011011;
		correct = 32'b01101100100100100111101010011110;
		#500; //1.4166577e+27 * -1.4044752e-32 = 1.4166577e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100101000001001010100110101011;
		x2 = 32'b01001001100010100110111000111101;
		correct = 32'b11100101000001001010100110101011;
		#500; //-3.9155137e+22 * 1134023.6 = -3.9155137e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011111100100111111110100011101;
		x2 = 32'b11101001111011100100011100000111;
		correct = 32'b11101001111011100100011100000111;
		#500; //6.267566e-20 * -3.600747e+25 = -3.600747e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001100001001011110111010011011;
		x2 = 32'b00000101011011100110010110110001;
		correct = 32'b00001100001001011111001001010101;
		#500; //1.278294e-31 * 1.1209384e-35 = 1.2784062e-31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111001000011111111110111111;
		x2 = 32'b01001101011101110011000100100101;
		correct = 32'b01001101011101110011000100100101;
		#500; //9.655893e-06 * 259199570.0 = 259199570.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101101101001010011101100101001;
		x2 = 32'b01010000100001111101000011001110;
		correct = 32'b01010000100001111101000011001110;
		#500; //-1.87846e-11 * 18228867000.0 = 18228867000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010010011101000010001001000010;
		x2 = 32'b10010100110010011100000010011111;
		correct = 32'b10010100110100010110000110110001;
		#500; //-7.703505e-28 * -2.0371789e-26 = -2.114214e-26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110110010010011000010100001;
		x2 = 32'b01010000100111111100011111101010;
		correct = 32'b01010000100111111100011111101010;
		#500; //7.567925e-35 * 21445431000.0 = 21445431000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000011110001011010100110000111;
		x2 = 32'b10011011110100000100110011111010;
		correct = 32'b01000011110001011010100110000111;
		#500; //395.32443 * -3.4460458e-22 = 395.32443
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111011000001111010010111100010;
		x2 = 32'b01110000010100101110111001010011;
		correct = 32'b01111011000001111010010111100101;
		#500; //7.043246e+35 * 2.6111987e+29 = 7.043248e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100110000001000011011011101;
		x2 = 32'b01001101110010110110110010100111;
		correct = 32'b11110100110000001000011011011101;
		#500; //-1.2202836e+32 * 426611940.0 = -1.2202836e+32
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100111011100101101001111111;
		x2 = 32'b01111001011111001000000010101111;
		correct = 32'b01111001011111001000000010101111;
		#500; //-1.5772912e-21 * 8.19418e+34 = 8.19418e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001111010011010011011010110100;
		x2 = 32'b00101000010111110010000110001001;
		correct = 32'b01001111010011010011011010110100;
		#500; //3442914300.0 * 1.23862585e-14 = 3442914300.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001010000110000101100111010;
		x2 = 32'b00100110101101010100011100000000;
		correct = 32'b00100110101101010100011100000000;
		#500; //-3.5823898e-38 * 1.2578643e-15 = 1.2578643e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001000101011111000000010011111;
		x2 = 32'b10101100101100101000100010010000;
		correct = 32'b10101100101100101000100010010000;
		#500; //1.0562668e-33 * -5.0742258e-12 = -5.0742258e-12
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001111110011001011000010101100;
		x2 = 32'b11100001011101000100101100011100;
		correct = 32'b11100001011101000100101100011100;
		#500; //6868261000.0 * -2.8165111e+20 = -2.8165111e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101100110010100010000001110011;
		x2 = 32'b11111000001001110100001010111101;
		correct = 32'b11111000001001110100001010111101;
		#500; //5.744788e-12 * -1.35698e+34 = -1.35698e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001111101001110010010010111111;
		x2 = 32'b11000011101010110110100001101011;
		correct = 32'b01001111101001110010010010111110;
		#500; //5608406500.0 * -342.81577 = 5608406000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000110001001110011000011100;
		x2 = 32'b01101101101010101011011001101000;
		correct = 32'b01101101101010101011011001101000;
		#500; //26427318000.0 * 6.604121e+27 = 6.604121e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101000110001100111001101011;
		x2 = 32'b11111101000000001001001100110000;
		correct = 32'b11111101000000001001001100110000;
		#500; //-1.3253836e-16 * -1.0681589e+37 = -1.0681589e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111011011110100011010000010;
		x2 = 32'b10011100101110010100101101101101;
		correct = 32'b11111111011011110100011010000010;
		#500; //-3.1805159e+38 * -1.226177e-21 = -3.1805159e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001010011001111110100001101111;
		x2 = 32'b00001111011110100001101110010000;
		correct = 32'b00001111011110100101010110001010;
		#500; //1.1165961e-32 * 1.233126e-29 = 1.2342426e-29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011001101010001100000110000111;
		x2 = 32'b01001000001110010011100100011100;
		correct = 32'b01001000001110010011100100011100;
		#500; //1.7448958e-23 * 189668.44 = 189668.44
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011000000010101000110001011011;
		x2 = 32'b11010101001010000101001100101011;
		correct = 32'b11011000000011010010110110101000;
		#500; //-609341700000000.0 * -11567197000000.0 = -620908900000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011010001010100101001101010100;
		x2 = 32'b11000011110110101100010010001010;
		correct = 32'b11000011110110101100010010001010;
		#500; //3.5222488e-23 * -437.53546 = -437.53546
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101110100101111100111010100001;
		x2 = 32'b01100010011110001001101101101000;
		correct = 32'b11101110100101111100111010100001;
		#500; //-2.3491018e+28 * 1.1464977e+21 = -2.3491018e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100000010000011110001100111;
		x2 = 32'b11101011111001000010110010101101;
		correct = 32'b11111100000010000011110001100111;
		#500; //-2.82951e+36 * -5.5169212e+26 = -2.82951e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100110001011101101001011111011;
		x2 = 32'b01011011001100010010111010010101;
		correct = 32'b11100110001011101101001011111000;
		#500; //-2.0639592e+23 * 4.987229e+16 = -2.0639586e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111100001000111101011110000100;
		x2 = 32'b11101011110000111111010010011000;
		correct = 32'b01111100001000111101011110000100;
		#500; //3.4028623e+36 * -4.737912e+26 = 3.4028623e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001111110010100111000100001100;
		x2 = 32'b11011100011110100001001010101000;
		correct = 32'b11011100011110100001001010101000;
		#500; //-1.9962282e-29 * -2.8155703e+17 = -2.8155703e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000000001001011011100010110100;
		x2 = 32'b01011000101000100000110101000011;
		correct = 32'b01011000101000100000110101000011;
		#500; //3.464172e-39 * 1425422700000000.0 = 1425422700000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001000101110011011010000100000;
		x2 = 32'b11011010001100011010110011001011;
		correct = 32'b11011010001100011010110011001011;
		#500; //1.117663e-33 * -1.2502765e+16 = -1.2502765e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011001000010100100000111101100;
		x2 = 32'b00110000100001000111111101110110;
		correct = 32'b11011001000010100100000111101100;
		#500; //-2432251800000000.0 * 9.640491e-10 = -2432251800000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001011111100010110110000010000;
		x2 = 32'b11001000110111110000001101000001;
		correct = 32'b11001011111101001110100000011101;
		#500; //-31643680.0 * -456730.03 = -32100410.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001111000010010110000100100110;
		x2 = 32'b01010010011110010111101011110100;
		correct = 32'b01010010011101110101010101101111;
		#500; //-2304845300.0 * 267877420000.0 = 265572560000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111010111110010011110110001;
		x2 = 32'b10000100000000001111111111110110;
		correct = 32'b00100111010111110010011110110001;
		#500; //3.0968984e-15 * -1.516386e-36 = 3.0968984e-15
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101010001000011001101001010001;
		x2 = 32'b10111101110101001100001100010011;
		correct = 32'b11101010001000011001101001010001;
		#500; //-4.884145e+25 * -0.1038877 = -4.884145e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101110111010000010001000001101;
		x2 = 32'b10100111011000111010101111010000;
		correct = 32'b00101110111010000010000001000110;
		#500; //1.0556187e-10 * -3.1595718e-15 = 1.05558715e-10
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000001101101001111010011000100;
		x2 = 32'b00010101000010110110110111010000;
		correct = 32'b00010101000010110110110111010000;
		#500; //6.647278e-38 * 2.8157453e-26 = 2.8157453e-26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100010011000001100011101101110;
		x2 = 32'b11001000110110101001111000000011;
		correct = 32'b01100010011000001100011101101110;
		#500; //1.0366103e+21 * -447728.1 = 1.0366103e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100011001111000010101011101100;
		x2 = 32'b10111101101010110100110100100110;
		correct = 32'b01100011001111000010101011101100;
		#500; //3.4710807e+21 * -0.08364324 = 3.4710807e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011001001001100100011100100001;
		x2 = 32'b11111000100100100101001100011011;
		correct = 32'b11111000100100100101001100011011;
		#500; //8.596363e-24 * -2.374253e+34 = -2.374253e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001000100011101001110100011010;
		x2 = 32'b00110000100010000111001011011111;
		correct = 32'b01001000100011101001110100011010;
		#500; //292072.8 * 9.927951e-10 = 292072.8
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010101110100100110011011001001;
		x2 = 32'b11101010101000000111101111001111;
		correct = 32'b11101010101000000111101111001111;
		#500; //-8.498049e-26 * -9.70064e+25 = -9.70064e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100100111101111001110101101011;
		x2 = 32'b10111010111101000011001110110101;
		correct = 32'b01100100111101111001110101101011;
		#500; //3.6541512e+22 * -0.0018631133 = 3.6541512e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100000101011110010011000100011;
		x2 = 32'b10010001010101100101010111000010;
		correct = 32'b11100000101011110010011000100011;
		#500; //-1.0096651e+20 * -1.690805e-28 = -1.0096651e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100101111111100111101001100;
		x2 = 32'b00101011000000001110011010001111;
		correct = 32'b11111100101111111100111101001100;
		#500; //-7.9674654e+36 * 4.57947e-13 = -7.9674654e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101101001100000100100110101100;
		x2 = 32'b10010000011001001010011100001001;
		correct = 32'b00101101001100000100100110101100;
		#500; //1.00208e-11 * -4.509375e-29 = 1.00208e-11
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101111000110101110011101011000;
		x2 = 32'b10011010110001001100010001010011;
		correct = 32'b11101111000110101110011101011000;
		#500; //-4.794037e+28 * -8.138088e-23 = -4.794037e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101111011111100011010100111;
		x2 = 32'b11100110001110111100000101110010;
		correct = 32'b11100110001110111100000101110010;
		#500; //1.7864703e-06 * -2.2166274e+23 = -2.2166274e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000100101000101001110011010000;
		x2 = 32'b01000010010001100111010111101001;
		correct = 32'b01000100101010001101000001111111;
		#500; //1300.9004 * 49.615147 = 1350.5155
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111100010100111111110110001000;
		x2 = 32'b01111000110111000000010000100110;
		correct = 32'b01111100010101011011010110010000;
		#500; //4.4028674e+36 * 3.569967e+34 = 4.438567e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000111000010000111000000011100;
		x2 = 32'b11110001110011001100111101001001;
		correct = 32'b11110001110011001100111101001001;
		#500; //34928.11 * -2.0283371e+30 = -2.0283371e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001001011011101000010010011;
		x2 = 32'b01101000010000010111110010001000;
		correct = 32'b01101000010000010111110010001000;
		#500; //3.8594626e-14 * 3.6548557e+24 = 3.6548557e+24
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101100110100100010111100001111;
		x2 = 32'b10001101011101011011110011001001;
		correct = 32'b01101100110100100010111100001111;
		#500; //2.0327732e+27 * -7.5723696e-31 = 2.0327732e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001010010111111110010000110100;
		x2 = 32'b00110111111001010101001011100001;
		correct = 32'b00110111111001010101001011100001;
		#500; //-1.077998e-32 * 2.733752e-05 = 2.733752e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001101000011101011101000001000;
		x2 = 32'b10001100010000111001101100001000;
		correct = 32'b11001101000011101011101000001000;
		#500; //-149659780.0 * -1.5068907e-31 = -149659780.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100111000011111110110101111001;
		x2 = 32'b01111001111110100011110110000100;
		correct = 32'b01111001111110100011110110000100;
		#500; //6.79679e+23 * 1.6241524e+35 = 1.6241524e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100011000111000010101010111111;
		x2 = 32'b11100000010011101001010100101001;
		correct = 32'b11100011000111110110010100010100;
		#500; //-2.8807723e+21 * -5.9543397e+19 = -2.9403158e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100000001110100100100000101111;
		x2 = 32'b01011101100010010001000110011000;
		correct = 32'b01100000001111101001000010111100;
		#500; //5.369212e+19 * 1.2346053e+18 = 5.492673e+19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001110100000000011001100000101;
		x2 = 32'b11011010000110110110101111000110;
		correct = 32'b11011010000110110110101111000110;
		#500; //-3.1603566e-30 * -1.093678e+16 = -1.093678e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111011000001010011011001011011;
		x2 = 32'b01111101011000010110000111100101;
		correct = 32'b01111101011000010110000111100101;
		#500; //-0.0020326588 * 1.8724037e+37 = 1.8724037e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100011000001000110111100000110;
		x2 = 32'b01101010101110001000010101011111;
		correct = 32'b01101010101110001000010101011111;
		#500; //-7.1792445e-18 * 1.1153609e+26 = 1.1153609e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011101100000000101001111110010;
		x2 = 32'b00001101100110001011011001001010;
		correct = 32'b00011101100000000101001111110010;
		#500; //3.3968115e-21 * 9.411608e-31 = 3.3968115e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100000000000100110101011000100;
		x2 = 32'b11101001111000010010100010010101;
		correct = 32'b11101001111000010010100010000101;
		#500; //3.7590156e+19 * -3.4024994e+25 = -3.4024957e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001111110111101010011111010010;
		x2 = 32'b10000111011111011101000010011001;
		correct = 32'b00001111110111101010011101010011;
		#500; //2.1955532e-29 * -1.9094906e-34 = 2.1955341e-29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011100100011110110000001010101;
		x2 = 32'b10100110010110000000110001110000;
		correct = 32'b11011100100011110110000001010101;
		#500; //-3.2285472e+17 * -7.495691e-16 = -3.2285472e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010110111011111111110001011110;
		x2 = 32'b10011111001111111000100001000010;
		correct = 32'b11010110111011111111110001011110;
		#500; //-131933590000000.0 * -4.0558533e-20 = -131933590000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111010100111111001100000100;
		x2 = 32'b10101010000001011100000001100111;
		correct = 32'b10110111010100111111001100000100;
		#500; //-1.26331615e-05 * -1.1879526e-13 = -1.26331615e-05
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001100111110101000100111100001;
		x2 = 32'b11100110111001101110000100110001;
		correct = 32'b11100110111001101110000100110001;
		#500; //-131354376.0 * -5.4514917e+23 = -5.4514917e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111101010011111010011110000000;
		x2 = 32'b01100101100100010000111010101100;
		correct = 32'b01100101100100010000111010101100;
		#500; //-0.05069685 * 8.562672e+22 = 8.562672e+22
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101011101101101100111001100;
		x2 = 32'b11010100110011110111000010000101;
		correct = 32'b11010100110011110111000010000101;
		#500; //1.16068674e-35 * -7127568000000.0 = -7127568000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111011010001110111010111001;
		x2 = 32'b01111000011101101011101001100000;
		correct = 32'b01111000011101101011101001100000;
		#500; //-1.6784556e+19 * 2.0016956e+34 = 2.0016956e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011111110011101000110001101;
		x2 = 32'b10011101010111000101001101000100;
		correct = 32'b10011101010111000101001101000100;
		#500; //-1.4683015e-36 * -2.9159805e-21 = -2.9159805e-21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000000111110100101100111110;
		x2 = 32'b00011111111100000110010110101000;
		correct = 32'b00011111111100000110010110101000;
		#500; //3.1415185e-29 * 1.0181213e-19 = 1.0181213e-19
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110111101011110100100000100;
		x2 = 32'b11110101100000011100010101111101;
		correct = 32'b11111110111101011110100100100100;
		#500; //-1.6343537e+38 * -3.290097e+32 = -1.634357e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011011110000010010000111101111;
		x2 = 32'b11100101111000011000011011010010;
		correct = 32'b11100101111000011000011011011110;
		#500; //-1.0872396e+17 * -1.3312743e+23 = -1.3312754e+23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110110000110010100110110011;
		x2 = 32'b11011010001111010000111110011001;
		correct = 32'b11011010001111010000111110011001;
		#500; //-5.8163073e-06 * -1.330398e+16 = -1.330398e+16
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100001101001100111101111000100;
		x2 = 32'b01101001111001011111001010111110;
		correct = 32'b01101001111001011111001010111110;
		#500; //1.1281358e-18 * 3.4748791e+25 = 3.4748791e+25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110100101100000110011101000;
		x2 = 32'b01100011011010110100010101100100;
		correct = 32'b11111110100101100000110011101000;
		#500; //-9.972561e+37 * 4.339985e+21 = -9.972561e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110001010100110010101111110101;
		x2 = 32'b01010100100110000111101010001110;
		correct = 32'b11110001010100110010101111110101;
		#500; //-1.04567165e+30 * 5239129000000.0 = -1.04567165e+30
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000100011110110101101000111011;
		x2 = 32'b01000111101000101000110000100110;
		correct = 32'b01000111101001001000001011011010;
		#500; //1005.40985 * 83224.3 = 84229.7
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010101011101111011101101001000;
		x2 = 32'b11100010011101110001000110110011;
		correct = 32'b11100010011101110001000110110011;
		#500; //17023984000000.0 * -1.1394053e+21 = -1.1394053e+21
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011110100111110000101100011100;
		x2 = 32'b11001100100100010111010111001011;
		correct = 32'b11001100100100010111010111001011;
		#500; //1.6839375e-20 * -76263000.0 = -76263000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101000101000001001100100011;
		x2 = 32'b11101110100000001010110011011000;
		correct = 32'b01111101000101000001001100100011;
		#500; //1.2301569e+37 * -1.9911518e+28 = 1.2301569e+37
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100110000001110000010011100;
		x2 = 32'b10011111000111111000001101011100;
		correct = 32'b00111100110000001110000010011100;
		#500; //0.023544602 * -3.3778218e-20 = 0.023544602
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110100101010000101001111010010;
		x2 = 32'b00100101000001101001110100000010;
		correct = 32'b00110100101010000101001111010010;
		#500; //3.1353426e-07 * 1.1675844e-16 = 3.1353426e-07
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011011101110000101101001010110;
		x2 = 32'b10100001111011000001001111010111;
		correct = 32'b11011011101110000101101001010110;
		#500; //-1.0378144e+17 * -1.5997234e-18 = -1.0378144e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000011000011111011010101000100;
		x2 = 32'b00100010011011001111000000000001;
		correct = 32'b00100010011011001111000000000001;
		#500; //4.2232006e-37 * 3.2111021e-18 = 3.2111021e-18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110110101100111000010101000000;
		x2 = 32'b10001000110100101001110000111001;
		correct = 32'b01110110101100111000010101000000;
		#500; //1.8205542e+33 * -1.2675643e-33 = 1.8205542e+33
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001001001111110100010010101110;
		x2 = 32'b00010111011001001001000101110001;
		correct = 32'b00010111011001001001000101110001;
		#500; //2.3023082e-33 * 7.3854346e-25 = 7.3854346e-25
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010010110001001010101010000110;
		x2 = 32'b01011000100010000100110111101011;
		correct = 32'b01011000100010000100000110100000;
		#500; //-422337250000.0 * 1198945900000000.0 = 1198523500000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011010111010110010101000101111;
		x2 = 32'b00010010010000000101001100010001;
		correct = 32'b00011010111010110010101010001111;
		#500; //9.7261873e-23 * 6.0686905e-28 = 9.726248e-23
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111000110011001001101101011111;
		x2 = 32'b11010110011101101010100101001000;
		correct = 32'b11010110011101101010100101001000;
		#500; //9.756418e-05 * -67801730000000.0 = -67801730000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011111101110100111101000101111;
		x2 = 32'b01100010001101001100010101110011;
		correct = 32'b01100010001110101001100101000100;
		#500; //2.6874208e+19 * 8.336604e+20 = 8.605346e+20
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001000010011100011010100010000;
		x2 = 32'b01010101111111110100001100111011;
		correct = 32'b01010101111111110100001100111011;
		#500; //211156.25 * 35083027000000.0 = 35083027000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001001111011100100110111111100;
		x2 = 32'b10110001010010000111101110110011;
		correct = 32'b01001001111011100100110111111100;
		#500; //1952191.5 * -2.9174145e-09 = 1952191.5
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100010100110000010101101000;
		x2 = 32'b11010100011101000110100101101111;
		correct = 32'b11010100111000111011011101101100;
		#500; //-3625315200000.0 * -4198963600000.0 = -7824279000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001001111101100011110111101111;
		x2 = 32'b00110011000110010100101001111110;
		correct = 32'b11001001111101100011110111101111;
		#500; //-2017213.9 * 3.569084e-08 = -2017213.9
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111000000000000100110000011;
		x2 = 32'b10101101011111011011011001010011;
		correct = 32'b11010111000000000000100110000011;
		#500; //-140778340000000.0 * -1.4421869e-11 = -140778340000000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011011010000001100000111011;
		x2 = 32'b00100010100000100100001010000110;
		correct = 32'b11111011011010000001100000111011;
		#500; //-1.2051043e+36 * 3.5307005e-18 = -1.2051043e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011001001100110011101111000100;
		x2 = 32'b11101110111111000001111001000100;
		correct = 32'b11101110111111000001111001000100;
		#500; //9.266153e-24 * -3.9013406e+28 = -3.9013406e+28
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011101000010011001010000110001;
		x2 = 32'b11101011011110110000110000110101;
		correct = 32'b11101011011110110000110000110101;
		#500; //-6.1960016e+17 * -3.0349803e+26 = -3.0349803e+26
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100100001101001001010000101;
		x2 = 32'b10100100110000001110000001010000;
		correct = 32'b10111100100001101001001010000101;
		#500; //-0.016427288 * -8.364673e-17 = -0.016427288
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011111110100010010010111000;
		x2 = 32'b11011100111100011011001111001101;
		correct = 32'b11011100111100011011001111001101;
		#500; //-1.470211e-36 * -5.442653e+17 = -5.442653e+17
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101111111110011101000000000111;
		x2 = 32'b11010110101010011011000000111110;
		correct = 32'b11101111111110011101000000000111;
		#500; //-1.5462651e+29 * -93287210000000.0 = -1.5462651e+29
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011110001110101100001011000011;
		x2 = 32'b00001011100101001101010111010000;
		correct = 32'b01011110001110101100001011000011;
		#500; //3.3643833e+18 * 5.7329236e-32 = 3.3643833e+18
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101100111011011010100110000111;
		x2 = 32'b11010101011110110000101001100100;
		correct = 32'b01101100111011011010100110000111;
		#500; //2.2985279e+27 * -17251378000000.0 = 2.2985279e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011001001100111011000110110;
		x2 = 32'b00101111111011000100001110110000;
		correct = 32'b11111011001001100111011000110110;
		#500; //-8.643189e+35 * 4.2976245e-10 = -8.643189e+35
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010110101001000100011100110010;
		x2 = 32'b11010001101011110001011101101100;
		correct = 32'b11010001101011110001011101101100;
		#500; //2.654056e-25 * -94001530000.0 = -94001530000.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100101011011110001101011101110;
		x2 = 32'b01001100111100011010100100101101;
		correct = 32'b01001100111100011010100100101101;
		#500; //2.073907e-16 * 126699880.0 = 126699880.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110110100111101001101110000;
		x2 = 32'b11101101011010001010100110001101;
		correct = 32'b11101101011010001010100110001101;
		#500; //7.968006e-35 * -4.5003435e+27 = -4.5003435e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100001101110100111111011001001;
		x2 = 32'b11111000000110100001000111011010;
		correct = 32'b11111000000110100001000111011010;
		#500; //1.263741e-18 * -1.2499622e+34 = -1.2499622e+34
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110011000011011010111110011011;
		x2 = 32'b11001100011010010000101100111000;
		correct = 32'b01110011000011011010111110011011;
		#500; //1.1225518e+31 * -61091040.0 = 1.1225518e+31
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100010111001101111111001100111;
		x2 = 32'b01111011111101011010000111111100;
		correct = 32'b01111011111101011010000111111100;
		#500; //6.2610984e-18 * 2.5507963e+36 = 2.5507963e+36
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110110011110111000010001010;
		x2 = 32'b00010111010010000101011010001100;
		correct = 32'b11111110110011110111000010001010;
		#500; //-1.3786727e+38 * 6.4732723e-25 = -1.3786727e+38
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111101100101001110010110111;
		x2 = 32'b00111001011000001001001110000010;
		correct = 32'b00111001011101101110011100011001;
		#500; //2.129223e-05 * 0.00021417256 = 0.00023546479
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101101101000100000111101110010;
		x2 = 32'b01101011001111010100101110001000;
		correct = 32'b01101101101001111111100111001110;
		#500; //6.2694055e+27 * 2.2884367e+26 = 6.498249e+27
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000011101111011110110110000;
		x2 = 32'b01001100101010101010000000110001;
		correct = 32'b01001100101010101010000000110001;
		#500; //4.885829e-29 * 89457030.0 = 89457030.0
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100100100110011110111001000;
		x2 = 32'b10101001110110101101100010001011;
		correct = 32'b10101001110110101101100010001011;
		#500; //-9.743614e-22 * -9.718709e-14 = -9.718709e-14
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001000011111011110000011101111;
		x2 = 32'b00110010101001010110000001010010;
		correct = 32'b01001000011111011110000011101111;
		#500; //259971.73 * 1.925233e-08 = 259971.73
					end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
		end
		end
		
endmodule