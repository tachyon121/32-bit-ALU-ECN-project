`timescale 1 ns/1 ps
    `include "alu.v"


    module div_tb ();
        reg clock;
        reg [31:0] X1, X2;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] x3;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .x1(X1),
                .x2(X2),
                .OpCode(op),
                .x3(x3)
            );
        /* create X1 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, X1, X2, op, x3);
            clock = 0;

    op = 3'b010;

		/* Display the operation */
		$display ("Opcode: 010, Operation: DIV");
		/* Test Cases!*/
		X1 = 32'b00100001110010011001000010000101;
		X2 = 32'b10100111001000101111000001010010;
		correct = 32'b10111010000111100101011111100011;
		#400; //1.3658544e-18 * -2.2612294e-15 = -0.0006040318
				
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00110111110001000010101110010010;
		X2 = 32'b00011011010011000111011100001011;
		correct = 32'b01011011111101011001110101001111;
		#400; //2.338531e-05 * 1.6912949e-22 = 1.3826866e+17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011001100011100001101000110000;
		X2 = 32'b11110000101011100010110001000110;
		correct = 32'b10101000010100001101110011001001;
		#400; //4999780000000000.0 * -4.3123132e+29 = -1.1594195e-14
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00010010011001100110101000111011;
		X2 = 32'b00010010100110111100001101011101;
		correct = 32'b00111111001111010101100010001110;
		#400; //7.2706142e-28 * 9.830036e-28 = 0.7396325
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10001001001000010001000101100001;
		X2 = 32'b10001101000111000001011010000111;
		correct = 32'b00111011100001000001010101110001;
		#400; //-1.9387842e-33 * -4.809833e-31 = 0.0040308763
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00110101001111010011011101010100;
		X2 = 32'b01010010101101011101100110100111;
		correct = 32'b00100010000001010010111101001000;
		#400; //7.04885e-07 * 390520340000.0 = 1.8049892e-18
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011100001111101001000101000001;
		X2 = 32'b01100111110011001001010010101010;
		correct = 32'b00110011111011100111011011101110;
		#400; //2.1455982e+17 * 1.9322103e+24 = 1.1104372e-07
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011110011000000000110010001101;
		X2 = 32'b10000101110010000011110001011110;
		correct = 32'b01011000000011110011100011110110;
		#400; //-1.1861057e-20 * -1.8830085e-35 = 629899200000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10110011111000111011101100010110;
		X2 = 32'b10010011010101100001111001010101;
		correct = 32'b01100000000010000010001100101111;
		#400; //-1.0604542e-07 * -2.7025552e-27 = 3.9238944e+19
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10001101100001001000100111001111;
		X2 = 32'b10001101001010111101010000100111;
		correct = 32'b00111111110001010111011010000101;
		#400; //-8.168304e-31 * -5.2948812e-31 = 1.5426794
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001111011000101011100000010100;
		X2 = 32'b01101011101111011010011110100010;
		correct = 32'b10100011000110010000001111011010;
		#400; //-3803714600.0 * 4.585572e+26 = -8.294962e-18
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010000001100111001101010100100;
		X2 = 32'b00111110110000101111101011011000;
		correct = 32'b11010000111010111100111111110000;
		#400; //-12053025000.0 * 0.38082004 = -31650185000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00100101100101011110011111110011;
		X2 = 32'b11100100001101101011000111101000;
		correct = 32'b10000000110100100000111000000111;
		#400; //2.6004555e-16 * -1.3480508e+22 = -1.9290486e-38
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11111000110011111100010000100001;
		X2 = 32'b11001101111101010101011111001011;
		correct = 32'b01101010010110001100101001111100;
		#400; //-3.3711982e+34 * -514521440.0 = 6.5521046e+25
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01111110001111101101100101100101;
		X2 = 32'b11010100101011111101000011110101;
		correct = 32'b11101001000010101111000111001010;
		#400; //6.3420524e+37 * -6041000000000.0 = -1.0498349e+25
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010100010111010100101111100001;
		X2 = 32'b10101100110010100101001111011110;
		correct = 32'b11100111000011000000000000011000;
		#400; //3801843200000.0 * -5.7504964e-12 = -6.6113304e+23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00001110100100101000010011101011;
		X2 = 32'b10110001000001010011110000010000;
		correct = 32'b10011101000011001100001100111101;
		#400; //3.6119774e-30 * -1.9388189e-09 = -1.8629782e-21
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11111110110100011101001110000001;
		X2 = 32'b01101110101110110110101010100100;
		correct = 32'b11001111100011110100111000011100;
		#400; //-1.3945342e+38 * 2.9001309e+28 = -4808521700.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011110011100001000101101001100;
		X2 = 32'b00111011001011010110110001101101;
		correct = 32'b10100010101100011000101001001010;
		#400; //-1.27343e-20 * 0.0026462332 = -4.8122365e-18
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001010110010001001100100010101;
		X2 = 32'b01101011100011011010001010101010;
		correct = 32'b00011110101101010100100101000011;
		#400; //6573194.5 * 3.424534e+26 = 1.919442e-20
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00001011011010011111110011100000;
		X2 = 32'b00101001011111111101010001111111;
		correct = 32'b00100001011010100010010010101010;
		#400; //4.506441e-32 * 5.6805685e-14 = 7.933081e-19
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01110011110101100010110100110011;
		X2 = 32'b11010010100001101110110010010011;
		correct = 32'b11100000110010110010111101110001;
		#400; //3.393763e+31 * -289747340000.0 = -1.1712836e+20
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100110001010000110100110010111;
		X2 = 32'b11011010010100111110100001010100;
		correct = 32'b11001011010010110111010001101001;
		#400; //1.9882634e+23 * -1.4911667e+16 = -13333609.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010100001111011101001111100010;
		X2 = 32'b01000101000001000000001111101101;
		correct = 32'b01001110101110000000110111001110;
		#400; //3261214500000.0 * 2112.2454 = 1543956200.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110101101010000111000000010011;
		X2 = 32'b01011011010010101000101100011101;
		correct = 32'b11011001110101001110010010011100;
		#400; //-4.2704053e+32 * 5.70109e+16 = -7490506700000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101010010100010010011001000001;
		X2 = 32'b10000011111000111111011101001100;
		correct = 32'b01100101111010101101111010010101;
		#400; //-1.8576201e-13 * -1.33986375e-36 = 1.3864246e+23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000110001000001000101111000111;
		X2 = 32'b01000101000111100011011010001000;
		correct = 32'b01000000100000011110001100110010;
		#400; //10274.944 * 2531.4082 = 4.058984
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011011110101111001000010110001;
		X2 = 32'b01101010101011100110100101101000;
		correct = 32'b00110000100111100011001111001100;
		#400; //1.2135242e+17 * 1.0542543e+26 = 1.1510735e-09
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010101000110000101100111100000;
		X2 = 32'b00100100010101001101010110011001;
		correct = 32'b01110000001101110011111111111001;
		#400; //10469486000000.0 * 4.6151096e-17 = 2.2685238e+29
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10000001011101111000011110001101;
		X2 = 32'b00000110101101001001000011001110;
		correct = 32'b10111010001011110111100000110110;
		#400; //-4.5463988e-38 * 6.7921246e-35 = -0.0006693633
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001010010110110001110011011110;
		X2 = 32'b10011100011011101111101011001101;
		correct = 32'b01101101011010101011011111011000;
		#400; //-3589943.5 * -7.9071747e-22 = 4.540109e+27
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000011100111110110100001110111;
		X2 = 32'b10100010101110001010110001110001;
		correct = 32'b11100000010111001111100111100110;
		#400; //318.81613 * -5.005588e-18 = -6.3692043e+19
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101011011011000110001110001100;
		X2 = 32'b10110100000000100111100011001110;
		correct = 32'b00110110111001111110100100001000;
		#400; //-8.398219e-13 * -1.2151142e-07 = 6.911465e-06
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10111001101001110000010010110011;
		X2 = 32'b00100001101000000000010111100001;
		correct = 32'b11010111100001011001100001110011;
		#400; //-0.00031856223 * 1.0843578e-18 = -293779620000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101110000011101110101111101111;
		X2 = 32'b10010100001010100010110000111011;
		correct = 32'b01011001010101110000000100101111;
		#400; //-3.2496613e-11 * -8.5915296e-27 = 3782401300000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10001111111000101101000110010100;
		X2 = 32'b10110111100001000111011101011010;
		correct = 32'b00010111110110110010101111011000;
		#400; //-2.2366047e-29 * -1.5791204e-05 = 1.4163611e-24
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11011100000101110010110011011110;
		X2 = 32'b00101100101111001011011010111000;
		correct = 32'b11101110110011010001001110111101;
		#400; //-1.7020821e+17 * 5.3635672e-12 = -3.1734145e+28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10100110001100011000100011001001;
		X2 = 32'b01000001100000110001101110111001;
		correct = 32'b10100100001011010101001101001011;
		#400; //-6.159459e-16 * 16.388536 = -3.7583947e-17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101010011000011010100001111001;
		X2 = 32'b00011010000100110110101111111110;
		correct = 32'b11001111110000111110110111011101;
		#400; //-2.0042465e-13 * 3.0486123e-23 = -6574291500.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11100111110110101000110100000000;
		X2 = 32'b01001010010101000111011011100010;
		correct = 32'b11011101000000111010101010110010;
		#400; //-2.0641538e+24 * 3481016.5 = -5.9297445e+17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01110110001111011110101011001100;
		X2 = 32'b01001110111010010100111110011000;
		correct = 32'b01100110110100000110001011100100;
		#400; //9.629945e+32 * 1957153800.0 = 4.9203822e+23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10001001100100011101010000010001;
		X2 = 32'b10000000000010100000000101100111;
		correct = 32'b01001010011010010011001010011011;
		#400; //-3.5106907e-33 * -9.18858e-40 = 3820710.8
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01101011101010011101100100011000;
		X2 = 32'b11010010101110000110010100001010;
		correct = 32'b11011000011010111100110111110011;
		#400; //4.1066732e+26 * -395984570000.0 = -1037079100000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101010000110001110011101100000;
		X2 = 32'b10011010011101100000000001001010;
		correct = 32'b11001111000111110001111001100010;
		#400; //1.3580586e-13 * -5.087184e-23 = -2669568500.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010110100111101010101010100000;
		X2 = 32'b01001111100111010101000111100010;
		correct = 32'b01000110100000010001100001111110;
		#400; //87227830000000.0 * 5278778400.0 = 16524.246
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101111010000000000010110111001;
		X2 = 32'b10001100110101110010110010001110;
		correct = 32'b01100001111001000111010010100101;
		#400; //-1.7464331e-10 * -3.315281e-31 = 5.2678285e+20
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11100000111110000110011110111110;
		X2 = 32'b01011101001010001101000111110000;
		correct = 32'b11000011001111000101011101111110;
		#400; //-1.4319587e+20 * 7.60298e+17 = -188.34177
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10111011111001110111111100011001;
		X2 = 32'b11110101011011010001101100000101;
		correct = 32'b00000101111110011111000110100111;
		#400; //-0.007064712 * -3.0056699e+32 = 2.3504617e-35
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00000110010100100110110011010010;
		X2 = 32'b00010010001010100001110110011011;
		correct = 32'b00110011100111100101010001111011;
		#400; //3.957656e-35 * 5.3679033e-28 = 7.372815e-08
					end  
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110000000000011100111100111000;
		X2 = 32'b01001100100110010000001000100110;
		correct = 32'b11100010110110010010111110000011;
		#400; //-1.6069631e+29 * 80220460.0 = -2.0031835e+21
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00100010100010100101111000010010;
		X2 = 32'b00010011000010010010101110000011;
		correct = 32'b01001111000000010001111000010001;
		#400; //3.7504576e-18 * 1.7313284e-27 = 2166231300.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00110101111010111000101111101011;
		X2 = 32'b01101100111010101010010001111110;
		correct = 32'b00001000100000000111111000111111;
		#400; //1.7549586e-06 * 2.2693235e+27 = 7.7334e-34
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01110000100101010011011100011000;
		X2 = 32'b10110011100110010101001110011000;
		correct = 32'b11111100011110010010001010110100;
		#400; //3.6943897e+29 * -7.139823e-08 = -5.174343e+36
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10000110111001100111001011011010;
		X2 = 32'b00011000100101100001101000111000;
		correct = 32'b10101101110001001000001111101101;
		#400; //-8.6685143e-35 * 3.8800565e-24 = -2.2341207e-11
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001111010111011101101101100111;
		X2 = 32'b11000000110111100011110111010101;
		correct = 32'b11001101111111111000111010011110;
		#400; //3722143500.0 * -6.945048 = -535942080.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010111111100110010100001011101;
		X2 = 32'b10011011001011001110110000000000;
		correct = 32'b11111100001100111111110101100111;
		#400; //534709370000000.0 * -1.4303762e-22 = -3.738243e+36
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101110010110001110111101001000;
		X2 = 32'b00001000011010001100101011100011;
		correct = 32'b11100101011011101000111110110000;
		#400; //-4.932524e-11 * 7.0053453e-34 = -7.041086e+22
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10110100011000100011000111111001;
		X2 = 32'b11100110111010001100010001000101;
		correct = 32'b00001100111110001100010111001001;
		#400; //-2.106607e-07 * -5.4960478e+23 = 3.8329488e-31
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10100110001111110000110010100110;
		X2 = 32'b01100011111011110100011111101111;
		correct = 32'b10000001110011000110010111111101;
		#400; //-6.628358e-16 * 8.8279104e+21 = -7.508411e-38
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011110110101100100100111010100;
		X2 = 32'b00100011010001000000101110110001;
		correct = 32'b00111011000010111110100100101101;
		#400; //2.2688666e-20 * 1.0627657e-17 = 0.00213487
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10010001000110101110011011111111;
		X2 = 32'b11000011001111000011100111111011;
		correct = 32'b00001101010100101010110101010001;
		#400; //-1.2219639e-28 * -188.22649 = 6.491987e-31
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10001111100000100100011001111101;
		X2 = 32'b11001000011101100001000010011010;
		correct = 32'b00000110100001111000100100001101;
		#400; //-1.2846141e-29 * -251970.4 = 5.0982734e-35
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101001000111101100010110110011;
		X2 = 32'b11001011111101101110011111010100;
		correct = 32'b10011100101001001001111011010100;
		#400; //3.5254524e-14 * -32362408.0 = -1.0893666e-21
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011001110010101011011000001100;
		X2 = 32'b10101100011101011100001101001000;
		correct = 32'b11101100110100110010011110101110;
		#400; //7132263500000000.0 * -3.4924997e-12 = -2.0421658e+27
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010000101111011011101111110001;
		X2 = 32'b01001111110110010010110110101001;
		correct = 32'b01000000010111111010011001100111;
		#400; //25465686000.0 * 7287296500.0 = 3.4945314
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100001110000001110010100001111;
		X2 = 32'b11110000100001110010010101110010;
		correct = 32'b10110000101101101011000111100010;
		#400; //4.4478503e+20 * -3.3460596e+29 = -1.32928e-09
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10111110001000010011110111011001;
		X2 = 32'b01101011101000010010101001111011;
		correct = 32'b10010010000000000000111101100010;
		#400; //-0.1574625 * 3.8967533e+26 = -4.040864e-28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101100110011001001011011100001;
		X2 = 32'b11010000010101110110010011100111;
		correct = 32'b00011011111100110010100010000111;
		#400; //-5.8147796e-12 * -14454857000.0 = 4.0227168e-22
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00110100101111111010010001000101;
		X2 = 32'b10000101111001000000011111000011;
		correct = 32'b11101110010101110010010111100100;
		#400; //3.5696044e-07 * -2.1443868e-35 = -1.6646271e+28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010111011110111010110011100101;
		X2 = 32'b00011000011011001101011010000100;
		correct = 32'b11111110100010000000010011011001;
		#400; //-276720000000000.0 * 3.0610588e-24 = -9.040009e+37
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000111100100111110101111110011;
		X2 = 32'b01100010111101011100101000000110;
		correct = 32'b00100100000110100001000100011010;
		#400; //75735.9 * 2.2670048e+21 = 3.3407912e-17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001011111001000100100011010001;
		X2 = 32'b10110000110110010100100110011111;
		correct = 32'b01011010100001100111101001100001;
		#400; //-29921698.0 * -1.5809752e-09 = 1.8926102e+16
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100000100010001101000110101000;
		X2 = 32'b11010001001010010100100000010011;
		correct = 32'b11001110110011101110100001100000;
		#400; //7.887077e+19 * -45441167000.0 = -1735667700.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010010010000010110100110000000;
		X2 = 32'b00101000110000100110010011001100;
		correct = 32'b01101000111111101011010100010000;
		#400; //207674670000.0 * 2.158204e-14 = 9.622569e+24
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00010010001010101001111000001110;
		X2 = 32'b00110110000100011110110110010100;
		correct = 32'b00011011100101011010011111111001;
		#400; //5.383736e-28 * 2.1744972e-06 = 2.4758532e-22
					end  
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10110000111100110011001011001001;
		X2 = 32'b00101001001101111011111110100001;
		correct = 32'b11000111001010010110100110111010;
		#400; //-1.7695011e-09 * 4.0800374e-14 = -43369.727
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100000101000110001000000010101;
		X2 = 32'b10100001110111101000111010111010;
		correct = 32'b11111110001110111001000010111011;
		#400; //9.399932e+19 * -1.5081085e-18 = -6.232928e+37
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011000110010000110011101010111;
		X2 = 32'b01011011000100101001001110111000;
		correct = 32'b00111101001011110000000100110101;
		#400; //1762769300000000.0 * 4.1257765e+16 = 0.04272576
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00001111011101111000110110011111;
		X2 = 32'b00010111110100010001110100011100;
		correct = 32'b00110111000101111000011101110011;
		#400; //1.22053155e-29 * 1.3513657e-24 = 9.031838e-06
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00110100001000000111000110001011;
		X2 = 32'b00110100111101111010101000000010;
		correct = 32'b00111110101001011101100000000000;
		#400; //1.4942468e-07 * 4.6131032e-07 = 0.32391357
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011011000111101010111011001101;
		X2 = 32'b00000010101011000100101001010100;
		correct = 32'b11010111111010111100011111110100;
		#400; //-1.3125935e-22 * 2.531579e-37 = -518488050000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10010000001011101100000010011001;
		X2 = 32'b10101001010001100101010010110110;
		correct = 32'b00100110011000011001000011000001;
		#400; //-3.446382e-29 * -4.4038307e-14 = 7.8258735e-16
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01101100010101111111001100101101;
		X2 = 32'b11011001000110101100010111011000;
		correct = 32'b11010010101100101001100000110110;
		#400; //1.0442697e+27 * -2722792400000000.0 = -383528930000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011011000010110011100110100111;
		X2 = 32'b10110110110100001011101001111000;
		correct = 32'b10100011101010101100000110010010;
		#400; //1.1516439e-22 * -6.220591e-06 = -1.8513417e-17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00001001101110011000100000001000;
		X2 = 32'b00001100100001111001111101011000;
		correct = 32'b00111100101011110001101010011000;
		#400; //4.4665053e-33 * 2.0895945e-31 = 0.021374986
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100000101000000101111110000011;
		X2 = 32'b01011000101101100101011010100010;
		correct = 32'b01000111011000010010100100111100;
		#400; //9.244879e+19 * 1603865600000000.0 = 57641.234
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100101111101111001011101010001;
		X2 = 32'b11101110100011100010111100011011;
		correct = 32'b10110110110111101110010001010001;
		#400; //1.4615198e+23 * -2.200191e+28 = -6.642695e-06
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010111001110010010001011001010;
		X2 = 32'b01011010101011110000000111111001;
		correct = 32'b10111100000001110110100001100000;
		#400; //-203559070000000.0 * 2.4630145e+16 = -0.008264631
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10001000000001110101001010100111;
		X2 = 32'b00111010110001101001100101000010;
		correct = 32'b10001100101011100110111101111011;
		#400; //-4.072224e-34 * 0.0015151876 = -2.687604e-31
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10010010101001001101011100001001;
		X2 = 32'b00011100010111011111010001011010;
		correct = 32'b10110101101111100001111111101101;
		#400; //-1.0402865e-27 * 7.3438583e-22 = -1.4165395e-06
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011000011000010110111011001011;
		X2 = 32'b10010011011011000010011010000100;
		correct = 32'b11000100011101000110000110101000;
		#400; //2.9136505e-24 * -2.9806377e-27 = -977.5259
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101110101111100101111111010101;
		X2 = 32'b00010011010110100101111111011111;
		correct = 32'b01011010110111110010110011101100;
		#400; //8.657223e-11 * 2.7562736e-27 = 3.1409156e+16
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10010000011000011000110000010000;
		X2 = 32'b01001011001010001110110001110000;
		correct = 32'b10000100101010101110011111100111;
		#400; //-4.4481326e-29 * 11070576.0 = -4.0179777e-36
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100111111101011101010010111010;
		X2 = 32'b00111000010010000001001100010100;
		correct = 32'b01101111000111010100010111110001;
		#400; //2.3218078e+24 * 4.7701484e-05 = 4.86737e+28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11100111100111110011101111000010;
		X2 = 32'b11110001000111011000011000110110;
		correct = 32'b00110110000000010110001110001010;
		#400; //-1.5039172e+24 * -7.8002236e+29 = 1.9280437e-06
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11100000100000111100101111011010;
		X2 = 32'b01000100101010011100110111110100;
		correct = 32'b11011011010001101011001010111110;
		#400; //-7.597539e+19 * 1358.436 = -5.5928575e+16
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10000101001101110110111011001100;
		X2 = 32'b00000100000110010000011100001111;
		correct = 32'b11000000100110010110111010110110;
		#400; //-8.624969e-36 * 1.7988305e-36 = -4.7947645
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001011100011001101010101001100;
		X2 = 32'b10111010000011011000001110001000;
		correct = 32'b11010000111111101100010011001111;
		#400; //18459288.0 * -0.0005398323 = -34194487000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001011010111110111011010110000;
		X2 = 32'b11100101001011100010011011001000;
		correct = 32'b00100101101001000011111001111001;
		#400; //-14644912.0 * -5.1400447e+22 = 2.8491798e-16
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101000101100001010111111101001;
		X2 = 32'b10100111101111001011001000010000;
		correct = 32'b01000000011011111011010101011010;
		#400; //-1.9616214e-14 * -5.237354e-15 = 3.7454438
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011101001010111101100110001111;
		X2 = 32'b01101001111101111010100111100111;
		correct = 32'b00110010101100011010001001100000;
		#400; //7.739429e+17 * 3.7425877e+25 = 2.0679352e-08
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000001000010101111111111000100;
		X2 = 32'b00011010110101110110011011110110;
		correct = 32'b11100101101001010011001001100101;
		#400; //-8.687443 * 8.908826e-23 = -9.751501e+22
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011111010010000001111010101011;
		X2 = 32'b10000111010011000110101111011010;
		correct = 32'b11010111011110101001110011111000;
		#400; //4.2377015e-20 * -1.5378949e-34 = -275552080000000.0
					end  
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011011111010110010011111011011;
		X2 = 32'b01111111011000111100110110111101;
		correct = 32'b00011100000001000010000110001010;
		#400; //1.3238088e+17 * 3.02803e+38 = 4.3718485e-22
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011100110011101010001100100100;
		X2 = 32'b11011010000011000101111001010000;
		correct = 32'b10000010001111000110110111111110;
		#400; //1.3674107e-21 * -9877549000000000.0 = -1.3843625e-37
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01101111000011001101100001100001;
		X2 = 32'b01011111000000101111100110010111;
		correct = 32'b01001111100010011010010101100101;
		#400; //4.3589487e+28 * 9.43774e+18 = 4618636000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101011110101101000000011100000;
		X2 = 32'b10100000001011100110010000110101;
		correct = 32'b11001011000111010111000100000010;
		#400; //1.5241385e-12 * -1.4771529e-19 = -10318082.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00110010100000010001000110110100;
		X2 = 32'b00111001000010001000100011011010;
		correct = 32'b00111000111100100000000010100001;
		#400; //1.5025627e-08 * 0.00013020952 = 0.000115395764
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01101110101000100011100110111001;
		X2 = 32'b11100001011001110100000011001110;
		correct = 32'b11001100101100111001010111100111;
		#400; //2.5103177e+28 * -2.6661672e+20 = -94154550.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01111010111011110101001111001100;
		X2 = 32'b11010011011111110001001000110100;
		correct = 32'b11100110111100000011001011101011;
		#400; //6.2132928e+35 * -1095522060000.0 = -5.671536e+23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110110010011110101000000010111;
		X2 = 32'b01110000011111011110110000001011;
		correct = 32'b11000101010100010000001001100111;
		#400; //-1.05120104e+33 * 3.1434026e+29 = -3344.1501
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11100111010100101101010111110101;
		X2 = 32'b01100001101010101110101101111100;
		correct = 32'b11000101000111011110010010000000;
		#400; //-9.956438e+23 * 3.9411437e+20 = -2526.2812
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10010101000111010110101010101101;
		X2 = 32'b00010111111110101101100111100000;
		correct = 32'b10111100101000001010010111010111;
		#400; //-3.179005e-26 * 1.6210871e-24 = -0.019610329
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10100110100101101110000010011110;
		X2 = 32'b01011111100101110101100100100011;
		correct = 32'b10000110011111110011010000100101;
		#400; //-1.0469223e-15 * 2.1811573e+19 = -4.799848e-35
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001110001011000010110000101011;
		X2 = 32'b01011000100011000101011100011111;
		correct = 32'b10110101000111010000100001111101;
		#400; //-722143940.0 * 1234446500000000.0 = -5.849941e-07
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00100100001100011110101110111011;
		X2 = 32'b00011011110100011110101011010001;
		correct = 32'b01000111110110001111101010111101;
		#400; //3.858043e-17 * 3.4727896e-22 = 111093.48
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101111101000010011010010110111;
		X2 = 32'b00001001110011101001011000111011;
		correct = 32'b01100101010001111100001110110110;
		#400; //2.9323186e-10 * 4.9733972e-33 = 5.8960072e+22
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100100010111100110010100111111;
		X2 = 32'b11001011110110000101001000001010;
		correct = 32'b11011000000000111001100000111101;
		#400; //1.6409891e+22 * -28353556.0 = -578759500000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110101101101000010000110011001;
		X2 = 32'b01110000111101001110011010011010;
		correct = 32'b11000100001111000100101110000110;
		#400; //-4.5668695e+32 * 6.0634498e+29 = -753.18005
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10110100001111010010010110010001;
		X2 = 32'b01010111110001011010111100101101;
		correct = 32'b10011011111101001111000110100110;
		#400; //-1.7615663e-07 * 434712330000000.0 = -4.0522576e-22
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00110010010111011110111001100010;
		X2 = 32'b10100001111101001110101111011011;
		correct = 32'b11001111111001111111100001001110;
		#400; //1.2918095e-08 * -1.6596514e-18 = -7783619600.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00001111000100100111000000110000;
		X2 = 32'b11000001110111110111011111010110;
		correct = 32'b10001100101001111100000110011110;
		#400; //7.219962e-30 * -27.933514 = -2.5846953e-31
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11101001110110100011000100010101;
		X2 = 32'b10101110010100111100000001001001;
		correct = 32'b01111011000000111110010010101100;
		#400; //-3.2972202e+25 * -4.814663e-11 = 6.848289e+35
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10111110001101011000101101101100;
		X2 = 32'b01110101101001101100000001111110;
		correct = 32'b10001000000010110101101011100000;
		#400; //-0.17728966 * 4.2276635e+32 = -4.1935614e-34
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010000110000101001101100101110;
		X2 = 32'b01110000101100011011100110011000;
		correct = 32'b10011111100011000010100001110111;
		#400; //-26119598000.0 * 4.4002573e+29 = -5.935925e-20
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001111011100111001011001101110;
		X2 = 32'b00010011101100100001011100011000;
		correct = 32'b11111011001011110001001101001101;
		#400; //-4086722000.0 * 4.495629e-27 = -9.090434e+35
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10110001111100010111101101101111;
		X2 = 32'b00100100010110101100001001001101;
		correct = 32'b11001101000011010100101110110111;
		#400; //-7.028056e-09 * 4.7435794e-17 = -148159340.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00000100011101100110010101001110;
		X2 = 32'b01000000101110111011001000010101;
		correct = 32'b00000011001010000000011111100100;
		#400; //2.8963678e-36 * 5.8654885 = 4.937982e-37
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010000001010101100101011010111;
		X2 = 32'b11011000011010001110101101111100;
		correct = 32'b00110111001110111011011101011011;
		#400; //-11461680000.0 * -1024392400000000.0 = 1.1188759e-05
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101100011101101111100001010010;
		X2 = 32'b10010101110110001111101110101001;
		correct = 32'b01010110000100011011000010000110;
		#400; //-3.5096548e-12 * -8.7638755e-26 = 40046837000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10100100010101001110010110110011;
		X2 = 32'b10000000000000100001101011101100;
		correct = 32'b01100110010010100100001100010000;
		#400; //-4.6164735e-17 * -1.93329e-40 = 2.3878878e+23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00000101010111100010111010010101;
		X2 = 32'b00100011010010010000010000011111;
		correct = 32'b00100001100011010111101001001001;
		#400; //1.04469456e-35 * 1.08971045e-17 = 9.5869e-19
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00000101111100010110011101001111;
		X2 = 32'b10000001110010101111101011101110;
		correct = 32'b11000011100110000011101011011011;
		#400; //2.270148e-35 * -7.456315e-38 = -304.4598
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11101000001101000000100000000110;
		X2 = 32'b01110010110011010010001001101010;
		correct = 32'b10110100111000001010110000011100;
		#400; //-3.400696e+24 * 8.126212e+30 = -4.1848477e-07
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000100001000100000000011011111;
		X2 = 32'b10100111101000100011001001100101;
		correct = 32'b11011011111111111011000111010110;
		#400; //648.0136 * -4.501867e-15 = -1.439433e+17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010000001000011000001111111110;
		X2 = 32'b11011001001010111110101011110100;
		correct = 32'b00110110011100001000001010100001;
		#400; //-10839128000.0 * -3024409700000000.0 = 3.5838823e-06
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10001110010101111000010001111000;
		X2 = 32'b00101011010011101100010011010110;
		correct = 32'b10100010100001010110101001110001;
		#400; //-2.6564577e-30 * 7.3459067e-13 = -3.616242e-18
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11100110101111011000101101100000;
		X2 = 32'b01001101100111101100110001000110;
		correct = 32'b11011000100110001100100010001100;
		#400; //-4.4754914e+23 * 333023420.0 = -1343896900000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000011101001001000111001000101;
		X2 = 32'b10011101001000010111111001111001;
		correct = 32'b01100110000000100110110100111101;
		#400; //-329.11148 * -2.1373557e-21 = 1.5398068e+23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10111001000101110000110101011101;
		X2 = 32'b10001010000101111001011101010011;
		correct = 32'b01101110011111110001011100000101;
		#400; //-0.0001440546 * -7.2988465e-33 = 1.9736627e+28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011000111001000011011001100101;
		X2 = 32'b11001001011110110010011111110101;
		correct = 32'b10001110111010001001110100101000;
		#400; //5.8991543e-24 * -1028735.3 = -5.734375e-30
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001101000101010110011001001000;
		X2 = 32'b11001101110111110100000010100111;
		correct = 32'b00111110101010110101000001100001;
		#400; //-156656770.0 * -468194530.0 = 0.33459762
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000001110010011111000110010001;
		X2 = 32'b10110010110111000000000001011010;
		correct = 32'b01001110011010101111110011001011;
		#400; //-25.242952 * -2.561153e-08 = 985608900.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11011000011010011101000011111100;
		X2 = 32'b11111101001110001010001001010011;
		correct = 32'b00011010101000100001100010100100;
		#400; //-1028335160000000.0 * -1.5338799e+37 = 6.704144e-23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100110011000000000110100011101;
		X2 = 32'b10110000001111011100011010111100;
		correct = 32'b11110101100101110001111000100001;
		#400; //2.64513e+23 * -6.904022e-10 = -3.8312886e+32
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11100111010111100000010011011110;
		X2 = 32'b11001001010110001111010000101100;
		correct = 32'b01011101100000101111110100001001;
		#400; //-1.04845514e+24 * -888642.75 = 1.1798388e+18
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01110011100010110001111000100010;
		X2 = 32'b01101000111000111010011111001011;
		correct = 32'b01001010000111000111000001010010;
		#400; //2.204408e+31 * 8.6005794e+24 = 2563092.5
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101000111110011000000100001100;
		X2 = 32'b00100010010110110101010100010100;
		correct = 32'b11000110000100011001101110100000;
		#400; //-2.7700518e-14 * 2.9725074e-18 = -9318.906
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10110000100001011100011100010001;
		X2 = 32'b00010111101011101011010001000011;
		correct = 32'b11011000010001000000011101101000;
		#400; //-9.733602e-10 * 1.1289991e-24 = -862144350000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011110001001100000110100011101;
		X2 = 32'b11000011110001101010111111001100;
		correct = 32'b10011001110101011111001101010010;
		#400; //8.7906786e-21 * -397.3734 = -2.212196e-23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000101001000011100100101001011;
		X2 = 32'b01001011011101001111000001110110;
		correct = 32'b00111001001010010001011110010010;
		#400; //2588.5808 * 16052342.0 = 0.00016125877
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000001001010111111001101000000;
		X2 = 32'b01010100111001010001011000110011;
		correct = 32'b00101011110000000010011010101010;
		#400; //10.746887 * 7871359600000.0 = 1.3653152e-12
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11100111001100101101100000101010;
		X2 = 32'b11010010000010100110001011000011;
		correct = 32'b01010100101001010110110000010110;
		#400; //-8.4456876e+23 * -148590610000.0 = 5683864000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001000101011011100000010010010;
		X2 = 32'b11110011100011111111001110001001;
		correct = 32'b10010100100110100111111110101001;
		#400; //355844.56 * -2.2809995e+31 = -1.5600379e-26
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01101011011010110000101010111101;
		X2 = 32'b11010001010000111101001011111001;
		correct = 32'b11011001100110011010001001111001;
		#400; //2.8414828e+26 * -52566135000.0 = -5405539000000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101110100101111101100001001111;
		X2 = 32'b00001110100101110111100110110100;
		correct = 32'b01011111100000000100111111110010;
		#400; //6.905109e-11 * 3.734157e-30 = 1.849175e+19
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11011010011000010110110110100000;
		X2 = 32'b01101100100000010101110001010000;
		correct = 32'b10101101010111110000111010100101;
		#400; //-1.5863101e+16 * 1.2510989e+27 = -1.2679334e-11
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010100001010110001000111011011;
		X2 = 32'b00101010100100110000110100000010;
		correct = 32'b11101001000101001110100001000000;
		#400; //-2938956000000.0 * 2.6121472e-13 = -1.1251112e+25
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011101000010100110010010101101;
		X2 = 32'b11000001010101101101011101101000;
		correct = 32'b10011011001001001110011111111010;
		#400; //1.8316196e-21 * -13.427589 = -1.3640718e-22
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10111101111100110110110010010011;
		X2 = 32'b00111101111011001111101110111111;
		correct = 32'b10111111100000110111101010010010;
		#400; //-0.11885943 * 0.11571454 = -1.027178
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10111111010011101010111001001000;
		X2 = 32'b01001101011010011111010100000101;
		correct = 32'b10110001011000100010011101011101;
		#400; //-0.8073468 * 245321810.0 = -3.2909704e-09
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000100011100100001100101000110;
		X2 = 32'b10110101000010111010110111100010;
		correct = 32'b01001110110111011101101100010001;
		#400; //-968.3949 * -5.203457e-07 = 1861060700.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000001110111110011010001101000;
		X2 = 32'b10110000000000101101101000101010;
		correct = 32'b01010001010110100101011011101001;
		#400; //-27.900589 * -4.7603754e-10 = 58610060000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11011101011000110101101110011110;
		X2 = 32'b00110000010110000110000010001000;
		correct = 32'b11101100100001100111111011101101;
		#400; //-1.02392886e+18 * 7.871752e-10 = -1.3007636e+27
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00111111101010010101100001010111;
		X2 = 32'b00000010111100101001001111011110;
		correct = 32'b01111100001100101011011100100001;
		#400; //1.3230084 * 3.5643576e-37 = 3.7117725e+36
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001001100110101100011100101000;
		X2 = 32'b01111110000100111001101101010010;
		correct = 32'b00001011000001100011011111111011;
		#400; //1267941.0 * 4.9050746e+37 = 2.5849576e-32
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010001110010100001010011000111;
		X2 = 32'b11010101001100000000101000001011;
		correct = 32'b10111100000100101110111101110100;
		#400; //108491500000.0 * -12097324000000.0 = -0.008968223
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10100010011111011000100001100001;
		X2 = 32'b00111011101010001101110111010100;
		correct = 32'b10100110010000000010110100110100;
		#400; //-3.4360092e-18 * 0.005153397 = -6.6674643e-16
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001000011100001110000110011100;
		X2 = 32'b10100011111110001011010001010100;
		correct = 32'b11100011111101111111001010001000;
		#400; //246662.44 * -2.6964586e-17 = -9.147644e+21
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010000110010111111001011000100;
		X2 = 32'b00100000001111001000110110111000;
		correct = 32'b01110000000010100111001101100011;
		#400; //27373478000.0 * 1.597111e-19 = 1.713937e+29
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101001011100100111110001000001;
		X2 = 32'b00011001011011001111111100010100;
		correct = 32'b01001111100000101111011011101101;
		#400; //5.3842567e-14 * 1.2252427e-23 = 4394441000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00111110011100110011010100011001;
		X2 = 32'b10000011000001101101100101011101;
		correct = 32'b11111010111001101101101011010001;
		#400; //0.23750724 * -3.962858e-37 = -5.993332e+35
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00111110001101110011001101011111;
		X2 = 32'b01110001000010101111110010000111;
		correct = 32'b00001100101010001011100000100000;
		#400; //0.1789069 * 6.882275e+29 = 2.5995315e-31
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110010001100101111000101110101;
		X2 = 32'b01101011110010001000010101101110;
		correct = 32'b11000101111001000111001110110010;
		#400; //-3.544335e+30 * 4.8483054e+26 = -7310.462
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10101000001100001000011110101010;
		X2 = 32'b00010000001100100110111001111010;
		correct = 32'b11010111011111010100010110001111;
		#400; //-9.79938e-15 * 3.5189418e-29 = -278475200000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00010100111001101010001000110001;
		X2 = 32'b01010011011011011110100100100101;
		correct = 32'b00000000111110000010101101100110;
		#400; //2.3288038e-26 * 1021818770000.0 = 2.2790771e-38
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011011001001100111011001011000;
		X2 = 32'b10010111100000001110010100110000;
		correct = 32'b11000011001001010100111001011100;
		#400; //1.3769437e-22 * -8.329661e-25 = -165.30609
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100100101111100010111010110100;
		X2 = 32'b10110101010100110100010001101100;
		correct = 32'b11101110111001100111001101100101;
		#400; //2.8065974e+22 * -7.870319e-07 = -3.5660528e+28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01101100101000011010010111101100;
		X2 = 32'b01001100110100100000111111011100;
		correct = 32'b01011111010001001111111110101000;
		#400; //1.5633648e+27 * 110132960.0 = 1.4195249e+19
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00010001110100001111100110011011;
		X2 = 32'b10100010110000010111000011010101;
		correct = 32'b10101110100010100100011101110000;
		#400; //3.2970445e-28 * -5.243222e-18 = -6.288203e-11
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000000010100110100100101101000;
		X2 = 32'b11011000101000011101000111011010;
		correct = 32'b00100111001001110010000011101011;
		#400; //-3.3013554 * -1423381400000000.0 = 2.319375e-15
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00001111011111000110001100000100;
		X2 = 32'b01000001110001101101000100110011;
		correct = 32'b00001101001000100111110100001111;
		#400; //1.2443629e-29 * 24.852148 = 5.007064e-31
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01110010001111001100000001111110;
		X2 = 32'b11111011010110010010101000010110;
		correct = 32'b10110110010111101000000110101011;
		#400; //3.738617e+30 * -1.127582e+36 = -3.3156055e-06
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110000011011011101000111101101;
		X2 = 32'b01010010000100110001111110110110;
		correct = 32'b11011101110011101110100000110011;
		#400; //-2.9440693e+29 * 157973050000.0 = -1.8636528e+18
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001101101100011000110111101001;
		X2 = 32'b11111111000001100011011011111010;
		correct = 32'b10001110001010010101010100110000;
		#400; //372358430.0 * -1.78402e+38 = -2.0871875e-30
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001100000001101010101010010110;
		X2 = 32'b10101110100111101001010011110011;
		correct = 32'b01011100110110010110010010011110;
		#400; //-35301976.0 * -7.211467e-11 = 4.895256e+17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011010011111111000001100010000;
		X2 = 32'b00011001000101100101000110100100;
		correct = 32'b11000000110110011001001100000101;
		#400; //-5.2838635e-23 * 7.7713054e-24 = -6.7991967
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11011111100000001100010110011101;
		X2 = 32'b10111011110111101101010101010001;
		correct = 32'b01100011000100111111000001000000;
		#400; //-1.855799e+19 * -0.0068003316 = 2.7289832e+21
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001001101000011100001011101111;
		X2 = 32'b00110001000011110000011100111111;
		correct = 32'b01011000000100001100001111001011;
		#400; //1325149.9 * 2.0813358e-09 = 636682400000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10001100001100000011001110010100;
		X2 = 32'b11001010000001111010010011110111;
		correct = 32'b00000001101001100100010101111101;
		#400; //-1.3574068e-31 * -2222397.8 = 6.107848e-38
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00010110001100110110111101010011;
		X2 = 32'b00111011000111110100101110100010;
		correct = 32'b00011010100100000010111011001100;
		#400; //1.4494633e-25 * 0.0024306555 = 5.963261e-23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010100001011011000011011000100;
		X2 = 32'b11010010010011110011011000101010;
		correct = 32'b01000001010101100110001000110100;
		#400; //-2981161300000.0 * -222491740000.0 = 13.398975
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01101011100111011100110111111011;
		X2 = 32'b10101111111000111101111001100111;
		correct = 32'b11111011001100010100100101000011;
		#400; //3.8154814e+26 * -4.1449086e-10 = -9.205225e+35
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011101010101100010010011011000;
		X2 = 32'b00000010111001000111100101111101;
		correct = 32'b11011001111011111111000101100000;
		#400; //-2.8341712e-21 * 3.357132e-37 = -8442239000000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010111101011101011101101011000;
		X2 = 32'b01010000101010111010001110010000;
		correct = 32'b01000110100000100100111001111001;
		#400; //384239320000000.0 * 23036985000.0 = 16679.236
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00010100111111100001101110100100;
		X2 = 32'b10100110011011000100111001010101;
		correct = 32'b10101110000010011010010010001111;
		#400; //2.5658348e-26 * -8.198511e-16 = -3.129635e-11
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110000001101111110101000100010;
		X2 = 32'b01001001111111111000001001111101;
		correct = 32'b11100101101110000100010001111010;
		#400; //-2.2767522e+29 * 2093135.6 = -1.08772325e+23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01010000001001111100000001110011;
		X2 = 32'b01010111011101111001101011001101;
		correct = 32'b00111000001011010111000010000111;
		#400; //11257630000.0 * 272244240000000.0 = 4.1351213e-05
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011100110011100111000001011010;
		X2 = 32'b11010000101110110000001101000001;
		correct = 32'b00001011100011010100101111010000;
		#400; //-1.3660979e-21 * -25100421000.0 = 5.4425294e-32
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01110011110100101110110111000101;
		X2 = 32'b11101001000010010011010010110010;
		correct = 32'b11001010010001001100011011001001;
		#400; //3.3423e+31 * -1.036698e+25 = -3223986.2
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00100100110111010101011111111010;
		X2 = 32'b00001000011000100001110111010000;
		correct = 32'b01011011111110101001100010110000;
		#400; //9.599251e-17 * 6.8044446e-34 = 1.4107325e+17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011101000101110101110110111010;
		X2 = 32'b11001010110001010011111001101000;
		correct = 32'b10010001110001000111010010111110;
		#400; //2.003314e-21 * -6463284.0 = -3.0995295e-28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001010110011011110000101011110;
		X2 = 32'b10011101100010010101001011000100;
		correct = 32'b01101100101111111110011100001001;
		#400; //-6746287.0 * -3.6349176e-21 = 1.8559669e+27
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110000000110000111000001100010;
		X2 = 32'b11111000001011000001100110000000;
		correct = 32'b00110111011000101100000100101111;
		#400; //-1.8871034e+29 * -1.3962379e+34 = 1.3515629e-05
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011110011100011101000000100100;
		X2 = 32'b00101011000010001101011100010110;
		correct = 32'b10110010111000100011000011111111;
		#400; //-1.2801476e-20 * 4.86154e-13 = -2.6332144e-08
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101110000101100100111110001110;
		X2 = 32'b00011000010011111111101001010001;
		correct = 32'b01010101001110010000010010000010;
		#400; //3.417671e-11 * 2.68805e-24 = 12714313000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011100111100011011011111101001;
		X2 = 32'b01011000101011010010000110100011;
		correct = 32'b00000011101100101011010100111100;
		#400; //1.5995582e-21 * 1522879800000000.0 = 1.0503509e-36
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001001001011110111011100000000;
		X2 = 32'b01010110111010101111010100100001;
		correct = 32'b00110001101111110010110111100010;
		#400; //718704.0 * 129169270000000.0 = 5.564048e-09
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10010100010101111111001111100101;
		X2 = 32'b10010100101010001010100100010100;
		correct = 32'b00111111001000111110010000011111;
		#400; //-1.0902826e-26 * -1.7030354e-26 = 0.6401996
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01101100010010100010111001000110;
		X2 = 32'b01001001110101110000100000110110;
		correct = 32'b01100001111100001011001101000011;
		#400; //9.7768614e+26 * 1761542.8 = 5.5501697e+20
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000101001010110000110110010011;
		X2 = 32'b01110110000010010000000110000111;
		correct = 32'b00001110100111111100111100011011;
		#400; //2736.8484 * 6.947028e+32 = 3.939596e-30
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11011001100111101111010100010101;
		X2 = 32'b11010111100000011010111111110100;
		correct = 32'b01000001100111001110001110100011;
		#400; //-5592814600000000.0 * -285185430000000.0 = 19.61115
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000011001010010111100010000000;
		X2 = 32'b00101001010101001010011110011010;
		correct = 32'b11011001010011000000001110001011;
		#400; //-169.4707 * 4.7218827e-14 = -3589049400000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10010010110111101111100011001110;
		X2 = 32'b10111111110101110011101011100000;
		correct = 32'b00010010100001001001101010101110;
		#400; //-1.4071505e-27 * -1.6814842 = 8.368503e-28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00111110111011100110110010000010;
		X2 = 32'b00011011100100001100110100101000;
		correct = 32'b01100010110100101100001001101000;
		#400; //0.4656716 * 2.395538e-22 = 1.9439124e+21
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000001111111011101101110011110;
		X2 = 32'b00010011111010110010111110101001;
		correct = 32'b11101101100010100010100101111101;
		#400; //-31.732235 * 5.9369337e-27 = -5.344886e+27
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01111011101111100110101010100011;
		X2 = 32'b01110110110100010111001001111101;
		correct = 32'b01000100011010001011110101001110;
		#400; //1.9773985e+36 * 2.1240472e+33 = 930.9579
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001000001111110001101011101111;
		X2 = 32'b01111011000111000100011111011001;
		correct = 32'b10001100100111001000010111001110;
		#400; //-195691.73 * 8.1145555e+35 = -2.4116136e-31
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011010011011110001100111000101;
		X2 = 32'b01010100001111000010011010001001;
		correct = 32'b00000101101000101010100101100101;
		#400; //4.9444858e-23 * 3232401500000.0 = 1.5296633e-35
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011110101101011110011001010001;
		X2 = 32'b01101101011001010010001100100101;
		correct = 32'b00110000110010110011100101111011;
		#400; //6.5536264e+18 * 4.4321596e+27 = 1.4786531e-09
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11000000010001110001111110111010;
		X2 = 32'b10001101101001011101001000111111;
		correct = 32'b01110010000110011011010011110011;
		#400; //-3.1113114 * -1.0219525e-30 = 3.0444775e+30
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10100101110010101010111011100011;
		X2 = 32'b00101001001010000111001000000111;
		correct = 32'b10111100000110100000010001010100;
		#400; //-3.5159922e-16 * 3.7402397e-14 = -0.009400446
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11001011000011010011001011001011;
		X2 = 32'b00110000110100011111011000000010;
		correct = 32'b11011001101011000010100011011011;
		#400; //-9253579.0 * 1.5276671e-09 = -6057327000000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010001000100011010111100000101;
		X2 = 32'b11100011110110101101111101110111;
		correct = 32'b00101100101010100110010101010010;
		#400; //-39106662000.0 * -8.074985e+21 = 4.8429394e-12
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011100100100000000011001100000;
		X2 = 32'b01000010100101100111001100010101;
		correct = 32'b10011001011101010001000101101100;
		#400; //-9.530769e-22 * 75.22477 = -1.26697214e-23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011010011001111111110111000100;
		X2 = 32'b01011010001001100111001110100111;
		correct = 32'b00111111101100100110011000111010;
		#400; //1.6324934e+16 * 1.1713002e+16 = 1.3937447
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11011111111001101110001011110011;
		X2 = 32'b00110110011110101100110100011111;
		correct = 32'b11101000111010111010110000100111;
		#400; //-3.3274254e+19 * 3.73723e-06 = -8.903454e+24
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10011001111001111001111100010111;
		X2 = 32'b00100011111110100010101100100101;
		correct = 32'b10110101011011010000010101000100;
		#400; //-2.3949096e-23 * 2.7123327e-17 = -8.829704e-07
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00111111100011110010000000000010;
		X2 = 32'b10101011100111110110101011110101;
		correct = 32'b11010011011001011101011000011100;
		#400; //1.1181643 * -1.1327316e-12 = -987139700000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10110101111010000000101001111000;
		X2 = 32'b00110010001101001111101010101100;
		correct = 32'b11000011001001000001110100110101;
		#400; //-1.7288394e-06 * 1.0534375e-08 = -164.11409
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00001010000010110011100011110000;
		X2 = 32'b00010110101100011000101010111110;
		correct = 32'b00110010110010001011111100011110;
		#400; //6.703315e-33 * 2.868345e-25 = 2.3369974e-08
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000101000011010110010111010110;
		X2 = 32'b00110000010011111001010111101000;
		correct = 32'b01010100001011100110000000100000;
		#400; //2262.3647 * 7.551919e-10 = 2995748000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01011001110110000011110111111001;
		X2 = 32'b00110101000110101100110001100001;
		correct = 32'b01100100001100101100111010000101;
		#400; //7608342000000000.0 * 5.766688e-07 = 1.3193607e+22
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01111011001011000001101110111110;
		X2 = 32'b01011110100111110111100111101011;
		correct = 32'b01011100000010100010001110001110;
		#400; //8.936377e+35 * 5.745737e+18 = 1.5553056e+17
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010010100101110000110111110000;
		X2 = 32'b11010110011111011110010101011000;
		correct = 32'b00111011100110000100111001101001;
		#400; //-324386950000.0 * -69790366000000.0 = 0.004648019
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b10110110010101011001010010000010;
		X2 = 32'b00111011011010110011001001011000;
		correct = 32'b10111010011010000111100010110001;
		#400; //-3.1825916e-06 * 0.0035888162 = -0.0008868082
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010111110111010010101000110001;
		X2 = 32'b10111100101000111110110110100101;
		correct = 32'b01011010101011001011000100100011;
		#400; //-486346560000000.0 * -0.020010779 = 2.430423e+16
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001010001001011111100110000101;
		X2 = 32'b11001111111000111110011100000010;
		correct = 32'b10111001101110100110111111111000;
		#400; //2719329.2 * -7647134700.0 = -0.00035560108
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11111011001001000111000101000010;
		X2 = 32'b01001110110001011001000110000101;
		correct = 32'b11101011110101010001001110101100;
		#400; //-8.538338e+35 * 1657324200.0 = -5.151882e+26
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11110010011000010000001010001001;
		X2 = 32'b11011001110011111101010010011011;
		correct = 32'b01011000000010101001010010100000;
		#400; //-4.4567803e+30 * -7312385300000000.0 = 609483800000000.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00111000000100110010100100001001;
		X2 = 32'b10010110000001000011101111001011;
		correct = 32'b11100001100011100111001011100111;
		#400; //3.5085748e-05 * -1.0681742e-25 = -3.2846466e+20
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00011010001010110101111000001010;
		X2 = 32'b10100100011010111011010000101001;
		correct = 32'b10110101001110100001111110100111;
		#400; //3.5437935e-23 * -5.1110104e-17 = -6.933646e-07
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00101011010001011011010101101000;
		X2 = 32'b01011000100100100011000101010110;
		correct = 32'b00010010001011010001101011100111;
		#400; //7.024021e-13 * 1285924800000000.0 = 5.4622334e-28
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01001001110011010100000111110011;
		X2 = 32'b10111011110101001101001111001111;
		correct = 32'b11001101011101101110010100001010;
		#400; //1681470.4 * -0.006494976 = -258887840.0
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b11010011111000011111111000100100;
		X2 = 32'b01111000110110011000111000110111;
		correct = 32'b10011010100001001111011011001110;
		#400; //-1941262800000.0 * 3.5300402e+34 = -5.4992655e-23
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b00110010101001100100100110000001;
		X2 = 32'b01001010000111110100001101000001;
		correct = 32'b00101000000001011010010101000011;
		#400; //1.935837e-08 * 2609360.2 = 7.4188185e-15
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01100011000110110011101101111111;
		X2 = 32'b11101010111111101110100010011000;
		correct = 32'b10110111100110111110010110100110;
		#400; //2.8635325e+21 * -1.5408278e+26 = -1.8584378e-05
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		X1 = 32'b01000101101100001001101011101001;
		X2 = 32'b10010001010100110110011101101010;
		correct = 32'b11110011110101011101110000111011;
		#400; //5651.364 * -1.6676832e-28 = -3.3887513e+31
					end 
 begin
			$display ("A      : %X2 %X2 %X2", X1[31], X1[30:23], X1[22:0]);
			$display ("B      : %X2 %X2 %X2", X2[31], X2[30:23], X2[22:0]);
			$display ("Output : %X2 %X2 %X2", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end
end
endmodule