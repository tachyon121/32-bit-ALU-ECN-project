`timescale 1 ps/1 ps
    `include "alu.v"


    module and_tb ();
        reg clk;
        reg [31:0] x1, x2;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] x3;
        wire [49:0] pro;

        alu U1 (
                .clk(clk),
                .x1(x1),
                .x2(x2),
                .OpCode(op),
                .x3(x3)
            );
        /* create x1 10Mhz clk */
        always
        #100 clk = ~clk; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clk, x1, x2, op, x3);
            clk = 0;

    op = 3'b100;

		/* Display the operation */
		$display ("Opcode: 100, Operation: AND");
		/* Test Cases!*/
		x1 = 32'b01110010110010001000000001010001;
		x2 = 32'b01001110001010001000000100001000;
		correct = 32'b01000010000010001000000000000000;
		
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110010111001001110000101000;
		x2 = 32'b00100011001111101110111011010000;
		correct = 32'b00100010000111001000110000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100101010101000110111010000000;
		x2 = 32'b11101101100001010101110100010000;
		correct = 32'b11100101000001000100110000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010010001100001000011000000;
		x2 = 32'b10011101001110011011000001000100;
		correct = 32'b10001000000000000001000001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100010101100100011110111101;
		x2 = 32'b00111001110100001010100100101101;
		correct = 32'b00010000010100000000000100101101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000001100011101110000111001;
		x2 = 32'b10100001010100010110011010011101;
		correct = 32'b00000000000100010100010000011001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100010101000111100100100000011;
		x2 = 32'b01111111110000110010111100011111;
		correct = 32'b01100010100000110000100100000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001001101101011111000010001010;
		x2 = 32'b00111011110101001011110000100111;
		correct = 32'b00001001100101001011000000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011110110110110111011100101100;
		x2 = 32'b10111010101001111001010011010000;
		correct = 32'b00011010100000110001010000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100000110010011100011100100;
		x2 = 32'b10110111010111011100100011101001;
		correct = 32'b10010100000110010000100011100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101001000110011001010011111;
		x2 = 32'b11100000011101001101101000010111;
		correct = 32'b01100000001000000001001000010111;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110110011110011000001100100000;
		x2 = 32'b11000110010011010010011101100101;
		correct = 32'b00000110010010010000001100100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100001001001011000110101111;
		x2 = 32'b10111011001100111010000000100011;
		correct = 32'b10010000001000001010000000100011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111001001101101100000000111;
		x2 = 32'b10001010101010001011100101111001;
		correct = 32'b10001010001000001001100000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001110010100000100001101101101;
		x2 = 32'b01000010110110010010100011011101;
		correct = 32'b01000010010100000000000001001101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101110100011111100011101101;
		x2 = 32'b01011110101111010011001000100011;
		correct = 32'b01011100100100010011000000100001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100011110110111000110110001100;
		x2 = 32'b01011011101100111011101010110101;
		correct = 32'b00000011100100111000100010000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101000001101010001011010101;
		x2 = 32'b10111110101100110010010011010101;
		correct = 32'b00111100000000100010000011010101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111010110110000111001000100;
		x2 = 32'b01100100100011100011011110100110;
		correct = 32'b01100100000010100000011000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000111100010000110000110101001;
		x2 = 32'b11010010100101000001101001001011;
		correct = 32'b01000010100000000000000000001001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110001000101110100010000000;
		x2 = 32'b00101010010101000000111101111101;
		correct = 32'b00101010000000000000100000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110101111100000100110001101;
		x2 = 32'b11001100010110101000010000011101;
		correct = 32'b00000100000110100000000000001101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110011100001001111010110100111;
		x2 = 32'b00010010110100111000110110111111;
		correct = 32'b00010010100000001000010110100111;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001101101110110110101001011001;
		x2 = 32'b11010110111111110101111111001101;
		correct = 32'b00000100101110110100101001001001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101011000000100001011100111001;
		x2 = 32'b11011101011110110010111100101001;
		correct = 32'b10001001000000100000011100101001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001101010100111011101011101110;
		x2 = 32'b01011100101101001011100101111001;
		correct = 32'b01001100000100001011100001101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100010110011000011101000000;
		x2 = 32'b00100010011001010001100110111100;
		correct = 32'b00100000010000010000000100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100101111100000110110000010;
		x2 = 32'b11000111110101000110100011101011;
		correct = 32'b11000100100101000000100010000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000000100111000111000111010;
		x2 = 32'b11100101101100011100110000100010;
		correct = 32'b11100000000100011000110000100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110001011100011010110000010110;
		x2 = 32'b10100000011001110111011011100010;
		correct = 32'b10100000011000010010010000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110011100000111000010001110;
		x2 = 32'b01100101001100001110000111111101;
		correct = 32'b00100100001100000110000010001100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000111000110101010011101010100;
		x2 = 32'b10011011011101111010000001110100;
		correct = 32'b00000011000100101010000001010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010010000001100010000110111111;
		x2 = 32'b00010111111001011110101110011011;
		correct = 32'b00010010000001000010000110011011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001111100110011000001101011101;
		x2 = 32'b01001000011101011011100001001010;
		correct = 32'b00001000000100011000000001001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011001100010110100101000000001;
		x2 = 32'b01010010000100000011001000110100;
		correct = 32'b01010000000000000000001000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101101101001001111101100010;
		x2 = 32'b00110010000000001000110110110110;
		correct = 32'b00110000000000001000110100100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011101011011100001010101010;
		x2 = 32'b00100000010000101001101101100101;
		correct = 32'b00100000000000001000001000100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011011101001000010011100000010;
		x2 = 32'b11000100010011000001101101110001;
		correct = 32'b11000000000001000000001100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110010111001110101001001010011;
		x2 = 32'b00000101101000011010111011010100;
		correct = 32'b00000000101000010000001001010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110011001000111101111110011110;
		x2 = 32'b01100111011100000111111111110000;
		correct = 32'b01100011001000000101111110010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100111011111010111000001111;
		x2 = 32'b10001001000110111100110010110100;
		correct = 32'b10000000000010111000110000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111110101100000011000101010010;
		x2 = 32'b00111001010100110100110011000011;
		correct = 32'b00111000000100000000000001000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100000001000100100011100100101;
		x2 = 32'b10100010111100001100001010011000;
		correct = 32'b10100000001000000100001000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111000010101110011000011001;
		x2 = 32'b01011100011011001111111110011000;
		correct = 32'b00010100000010001110011000011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000000100001110010011010110101;
		x2 = 32'b00010110101101001010010001001000;
		correct = 32'b00000000100001000010010000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100110110010011000110000011010;
		x2 = 32'b10011001010100000010000111011101;
		correct = 32'b10000000010000000000000000011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111111101101111111101001001100;
		x2 = 32'b11000000111000011000101001111011;
		correct = 32'b00000000101000011000101001001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100100111110100001110101100100;
		x2 = 32'b10101011011101000011110111111001;
		correct = 32'b00100000011100000001110101100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000101000000001101101110101011;
		x2 = 32'b00001101101101101011110110110111;
		correct = 32'b00000101000000001001100110100011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111110100101010110010000101;
		x2 = 32'b10110110100111001010010110101101;
		correct = 32'b10110110100100001010010010000101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011100100010011110101111100101;
		x2 = 32'b10000100010101101101001000011000;
		correct = 32'b00000100000000001100001000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111011011001000100100000000101;
		x2 = 32'b00101101101111110100011110000000;
		correct = 32'b00101001001001000100000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011001110010111011000110000110;
		x2 = 32'b11000100111110111101010100001010;
		correct = 32'b01000000110010111001000100000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001011101010001100110010000011;
		x2 = 32'b00100110101100011000010000010010;
		correct = 32'b00000010101000001000010000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010111001110010010000010111111;
		x2 = 32'b11101001010000001011101100110010;
		correct = 32'b01000001000000000010000000110010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000010110110010010010000111001;
		x2 = 32'b11000100111000111010111010000101;
		correct = 32'b00000000110000010010010000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101000100101010101110101110;
		x2 = 32'b01010001100010111110001001000100;
		correct = 32'b01010001000000101010001000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110100001010100011011111101000;
		x2 = 32'b00011101100111000111111111000011;
		correct = 32'b00010100000010000011011111000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001010100011110110000111101;
		x2 = 32'b01111011000011100001000101100111;
		correct = 32'b01100001000000000000000000100101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011010011010111001011110111111;
		x2 = 32'b10001110000000110101010011010101;
		correct = 32'b10001010000000110001010010010101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000100100110001011110111111111;
		x2 = 32'b00011010001100011111101001000001;
		correct = 32'b00000000000100001011100001000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111011111000010011000011101101;
		x2 = 32'b00111001011111111011111111100010;
		correct = 32'b00111001011000010011000011100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001011110101010101100001111011;
		x2 = 32'b01101111110010000000111000010011;
		correct = 32'b01001011110000000000100000010011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010011001001011111001000101000;
		x2 = 32'b01100111011101101110010101111011;
		correct = 32'b01000011001001001110000000101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101111000101111010100101001111;
		x2 = 32'b10000000011100110100101010100100;
		correct = 32'b00000000000100110000100000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111010011100111001000001000111;
		x2 = 32'b01010010100000101011000100000010;
		correct = 32'b01010010000000101001000000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000001111010101101100100000101;
		x2 = 32'b01010100101011101011101100010001;
		correct = 32'b00000000101010101001100100000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000000111100101011111001010110;
		x2 = 32'b11000111010001100100000110010001;
		correct = 32'b00000000010000100000000000010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111010001001111101110011110000;
		x2 = 32'b11110001100101100111111111000010;
		correct = 32'b01110000000001100101110011000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011101110000010110000110111100;
		x2 = 32'b10001110000100011010001101011010;
		correct = 32'b00001100000000010010000100011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101001111100101000000010000;
		x2 = 32'b11110101010011111101111101001111;
		correct = 32'b00110101000011100101000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110000111011000001000111010;
		x2 = 32'b01000110110101001010011110100111;
		correct = 32'b00000110000101001000001000100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111001101001110000000010110;
		x2 = 32'b00001001000110110010111110011011;
		correct = 32'b00000001000100000010000000010010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000101011000110100011000100000;
		x2 = 32'b01001001111001010111000001100100;
		correct = 32'b01000001011000010100000000100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100110100011101110101111110;
		x2 = 32'b00001111110001100100101010011000;
		correct = 32'b00000100110000000100100000011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010011000111101010101010011;
		x2 = 32'b11010001001111100101110100110110;
		correct = 32'b10000000001000100101010100010010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101110101110010101100100110110;
		x2 = 32'b10000110001001100011001101111000;
		correct = 32'b00000110001000000001000100110000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010010011000011011101001000101;
		x2 = 32'b01000001101110100110000101110011;
		correct = 32'b00000000001000000010000001000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001100101100010101000100000111;
		x2 = 32'b11011100000011001111100010000001;
		correct = 32'b11001100000000000101000000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100000000001100000000000001100;
		x2 = 32'b00001111111101011100110111011101;
		correct = 32'b00000000000001000000000000001100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001101011011011010111010111;
		x2 = 32'b11010111100101110001000110101100;
		correct = 32'b00000001100001010001000110000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111011011100011000011000101110;
		x2 = 32'b10100000010000001000010000000010;
		correct = 32'b00100000010000001000010000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101111110101010010000110111;
		x2 = 32'b10111010011110000110111011001111;
		correct = 32'b10100000011110000010010000000111;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111111100001001000001101110;
		x2 = 32'b10000110001001000001010010111101;
		correct = 32'b10000110001000000001000000101100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010000011001011110111010110;
		x2 = 32'b11000101001001011000001111001101;
		correct = 32'b01000000000001001000000111000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110110010001111010100100010010;
		x2 = 32'b10110100001111011111100100000100;
		correct = 32'b00110100000001011010100100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000000000001011100100110101;
		x2 = 32'b00011110011000001000001000100011;
		correct = 32'b00011000000000001000000000100001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011101010011000000001110101101;
		x2 = 32'b10010011010000100000110011001011;
		correct = 32'b00010001010000000000000010001001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101000101110100101001111101101;
		x2 = 32'b00111111110110110100011101111111;
		correct = 32'b00101000100110100100001101101101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100111010010000001011001110;
		x2 = 32'b10111111100101000111000100110000;
		correct = 32'b10011100100000000000000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101111000111011100001100001100;
		x2 = 32'b01100110111011100001110010001001;
		correct = 32'b01100110000011000000000000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100011100100010101100100010101;
		x2 = 32'b11110101101100001100001000010010;
		correct = 32'b01100001100100000100000000010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001001111011001110011001011011;
		x2 = 32'b01011110001010001111111100000111;
		correct = 32'b00001000001010001110011000000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101100110011010101101110111;
		x2 = 32'b01011100010000010011111111100010;
		correct = 32'b01010100000000010010101101100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111110110001001100010001001001;
		x2 = 32'b00101101001111110110001110010110;
		correct = 32'b00101100000001000100000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010000111100000110000001110100;
		x2 = 32'b10011000001001000001100010011111;
		correct = 32'b10010000001000000000000000010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001111110001101001000011111;
		x2 = 32'b01000101010100110010111100110001;
		correct = 32'b01000001010100000000001000010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111111011100010110001110011111;
		x2 = 32'b01110100110111011110101011000110;
		correct = 32'b00110100010100010110001010000110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110000000001011001011010110010;
		x2 = 32'b11011100001001110011010111000101;
		correct = 32'b00010000000001010001010010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110100100001100110010011011;
		x2 = 32'b11000000000110011010111110010111;
		correct = 32'b10000000000100001000110010010011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000111010111011110111010010011;
		x2 = 32'b01010000011011010111101000110011;
		correct = 32'b01000000010011010110101000010011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011011011011111100010001110001;
		x2 = 32'b01000010000001101101100100010011;
		correct = 32'b01000010000001101100000000010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010100001011110011010110010010;
		x2 = 32'b01101111110000100100001010110001;
		correct = 32'b00000100000000100000000010010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010111100101101011100101001101;
		x2 = 32'b10100110011010111010100101100001;
		correct = 32'b00000110000000101010100101000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001000110110011010011000011100;
		x2 = 32'b01011111010001000110111100110101;
		correct = 32'b00001000010000000010011000010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011101001011100010000110101;
		x2 = 32'b10001100001001011001110010110101;
		correct = 32'b00001000001001011000010000110101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010111011100101111100101101101;
		x2 = 32'b01100111110000001100011110100000;
		correct = 32'b00000111010000001100000100100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010010011100001000010000001101;
		x2 = 32'b01111101111101101100001000110010;
		correct = 32'b00010000011100001000000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010001101011101101000010010001;
		x2 = 32'b01000111011001011010110000110101;
		correct = 32'b00000001001001001000000000010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000100110111011100010000100000;
		x2 = 32'b11110101001011101011001001100001;
		correct = 32'b01000100000011001000000000100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110001111110000101110111011111;
		x2 = 32'b00111011001101100111111111100010;
		correct = 32'b00110001001100000101110111000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011101110011100000011100101010;
		x2 = 32'b10100010000011100100101001001001;
		correct = 32'b10000000000011100000001000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100001111000111100111111110000;
		x2 = 32'b00011010011101011101011010001111;
		correct = 32'b00000000011000011100011010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100011111110011111111101000;
		x2 = 32'b01100100000000011101011001111100;
		correct = 32'b01000100000000010001011001101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100101100010010001001010111;
		x2 = 32'b10001010001110101110010001110010;
		correct = 32'b10000000001100000010000001010010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111011100100000001110110000;
		x2 = 32'b10010111010000111010100101010011;
		correct = 32'b10010111010000100000000100010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111000010100101011000001101010;
		x2 = 32'b11000000010110101100001000100101;
		correct = 32'b01000000010100101000000000100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000000101111111001000101011;
		x2 = 32'b00001111001001100011000100000111;
		correct = 32'b00000000000001100011000000000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010111001001000100110001111111;
		x2 = 32'b10001100010100110110101111111101;
		correct = 32'b00000100000000000100100001111101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000110010010000000110110100100;
		x2 = 32'b01010110000001110101101111100111;
		correct = 32'b00000110000000000000100110100100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011111010111010000110110110010;
		x2 = 32'b00001110001001110000111101001011;
		correct = 32'b00001110000001010000110100000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010101101100110101100111001010;
		x2 = 32'b10010110110010100010001111100101;
		correct = 32'b10010100100000100000000111000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101001101101000000010101110101;
		x2 = 32'b01111110010110110000010110100101;
		correct = 32'b01101000000100000000010100100101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100000010010101110011010110110;
		x2 = 32'b11010001110010101010100110010111;
		correct = 32'b01000000010010101010000010010110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101011101001101101100000101000;
		x2 = 32'b00001011000001101011000110010100;
		correct = 32'b00001011000001101001000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011110000011110001100000011011;
		x2 = 32'b10110001110011011101111101110010;
		correct = 32'b10010000000011010001100000010010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001100110010011010011110010110;
		x2 = 32'b01001011000010001010110011110110;
		correct = 32'b00001000000010001010010010010110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011111001111001110011001000;
		x2 = 32'b00110000110000111011011101000011;
		correct = 32'b00000000110000111001010001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001011011100101000010000111;
		x2 = 32'b10110101100010001111100111100101;
		correct = 32'b10000001000010000101000010000101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110010001111001000111000100110;
		x2 = 32'b11110011000011010110101101110000;
		correct = 32'b10110010000011000000101000100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101100110111101110101010101100;
		x2 = 32'b10011100110110010110100010011010;
		correct = 32'b10001100110110000110100010001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000111010100011111010110111110;
		x2 = 32'b01000011111111000100110111101110;
		correct = 32'b00000011010100000100010110101110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110110001111101011010011000110;
		x2 = 32'b01101011000011110100101000110011;
		correct = 32'b00100010000011100000000000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101110101111101001110101001000;
		x2 = 32'b01100101000100000011110000101110;
		correct = 32'b00100100000100000001110000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011101011000011001010100000111;
		x2 = 32'b01010110101011100011111100100001;
		correct = 32'b00010100001000000001010100000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011001101101011111010110010100;
		x2 = 32'b10001111011010100000100101000100;
		correct = 32'b00001001001000000000000100000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101101010100110110101010110;
		x2 = 32'b00110100000101001000100000010000;
		correct = 32'b00110100000000000000100000010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101110100010001101011000011100;
		x2 = 32'b01010001011011101001001110010010;
		correct = 32'b01000000000010001001001000010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100110001001101010101110011101;
		x2 = 32'b00011011011000110001111110000111;
		correct = 32'b00000010001000100000101110000101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111110001010111001011000001;
		x2 = 32'b10000101100000100011111100001110;
		correct = 32'b10000101100000000011001000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100011111111111000111010000;
		x2 = 32'b11001000010101000000100110000011;
		correct = 32'b10001000010101000000000110000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101001100011000101110111010;
		x2 = 32'b11111001111100001000101010001100;
		correct = 32'b01110001001100001000101010001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110000011100001000111011011;
		x2 = 32'b00001000001111000110110101000000;
		correct = 32'b00000000000011000000000101000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001010010111101101010111110111;
		x2 = 32'b00011111101011001010100001000000;
		correct = 32'b00001010000011001000000001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011011101000111001101101101;
		x2 = 32'b00111010000111010101101101111100;
		correct = 32'b00100010000101000101001101101100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101010110111100011100110010011;
		x2 = 32'b00000111100111110000100101010000;
		correct = 32'b00000010100111100000100100010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101001010101101100100011010;
		x2 = 32'b01010111010000100101110100110001;
		correct = 32'b01010101000000100101100100010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101101001101101011010101101111;
		x2 = 32'b00001011111110000010101101010110;
		correct = 32'b00001001001100000010000101000110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011100010000000000010110111100;
		x2 = 32'b10010010011000100100111011010111;
		correct = 32'b00010000010000000000010010010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110101011110001111100101011101;
		x2 = 32'b01001111001010000110100111010011;
		correct = 32'b00000101001010000110100101010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110000010101111101011011110;
		x2 = 32'b01010111101001111111011100110010;
		correct = 32'b01010110000000101111001000010010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001101010110111001010110001110;
		x2 = 32'b00010011001010011011001010101001;
		correct = 32'b00000001000010011001000010001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000011010110001101001001111010;
		x2 = 32'b00110100110001110010011001010101;
		correct = 32'b00000000010000000000001001010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111011100011110000011011001111;
		x2 = 32'b11001110101010110000111011110001;
		correct = 32'b01001010100010110000011011000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010001001000101111000101011101;
		x2 = 32'b10101111110000001110001010000001;
		correct = 32'b00000001000000001110000000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110100101011101101101010110000;
		x2 = 32'b11100001010111110011010101111000;
		correct = 32'b10100000000011100001000000110000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111010000011110011100100101110;
		x2 = 32'b01000010001111110000011110010000;
		correct = 32'b01000010000011110000000100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011111111110000111110010011;
		x2 = 32'b01110110100111000110010000101001;
		correct = 32'b01100010100111000000010000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100110000100011011110101000;
		x2 = 32'b10110111101000001100010011111101;
		correct = 32'b10010100100000000000010010101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111100111110011101100101011;
		x2 = 32'b00000111100001110011100010011100;
		correct = 32'b00000111100001110011100000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111001011011000001001001001001;
		x2 = 32'b10001000101111001000010011000100;
		correct = 32'b10001000001011000000000001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101010101111111101001110100101;
		x2 = 32'b10111011110010100101111001010100;
		correct = 32'b10101010100010100101001000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010110100101001011110001100111;
		x2 = 32'b00010000100110100111101110110101;
		correct = 32'b00010000100100000011100000100101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110111110101110100010001000100;
		x2 = 32'b00111011011010110011010011100010;
		correct = 32'b00110011010000110000010001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001001101001010011111100010001;
		x2 = 32'b10010110010111011111001111111010;
		correct = 32'b00000000000001010011001100010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010001111010011111111100101011;
		x2 = 32'b11111000110110101001001011101110;
		correct = 32'b00010000110010001001001000101010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000101011100011001110000001000;
		x2 = 32'b11100111001001111000110111000100;
		correct = 32'b10000101001000011000110000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000011001011001110000111001011;
		x2 = 32'b01000001101100110101110111000000;
		correct = 32'b01000001001000000100000111000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011101011100010100011101010111;
		x2 = 32'b01001011100111010000011110011010;
		correct = 32'b00001001000100010000011100010010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101001000000000010001111111110;
		x2 = 32'b11111010010110010110011011001110;
		correct = 32'b11101000000000000010001011001110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101111110100110100111000001110;
		x2 = 32'b11101010111001111110011111001001;
		correct = 32'b01101010110000110100011000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001011110011100001010010010000;
		x2 = 32'b01101101011100111001110111001101;
		correct = 32'b00001001010000100001010010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010011100000100100101101100101;
		x2 = 32'b00100010100010011000000000011001;
		correct = 32'b00000010100000000000000000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100111101011011111011011000111;
		x2 = 32'b11000110000100110001100001100011;
		correct = 32'b10000110000000010001000001000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010101111100011010011100010;
		x2 = 32'b01011011000101010101001100100011;
		correct = 32'b01000010000101000001000000100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110100011010010111101110000110;
		x2 = 32'b01100110111111110001001001011011;
		correct = 32'b00100100011010010001001000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010111110011001011010101101110;
		x2 = 32'b01111010101001000000100010010011;
		correct = 32'b00010010100001000000000000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001101110100100101000010010111;
		x2 = 32'b10011100101000100000101100110111;
		correct = 32'b00001100100000100000000000010111;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010110111011011010110011000100;
		x2 = 32'b01100010111100011110110010101011;
		correct = 32'b00000010111000011010110010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101011111001100101010010000001;
		x2 = 32'b00001110100110000010000110100010;
		correct = 32'b00001010100000000000000010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101111011000001100111010001011;
		x2 = 32'b01110011011110001100000001001000;
		correct = 32'b01100011011000001100000000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111111010110100100110000110;
		x2 = 32'b01001001000000001001101001100100;
		correct = 32'b01001001000000000000100000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110001100101110010100101000101;
		x2 = 32'b11011001110110001110011110011000;
		correct = 32'b00010001100100000010000100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001010111011010001011011101101;
		x2 = 32'b01011000101101101101001001101101;
		correct = 32'b01001000101001000001001001101101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011110101101111110110000000;
		x2 = 32'b11111100101010000110110001010100;
		correct = 32'b01001000100000000110110000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011001100110101000000101000011;
		x2 = 32'b00011001101011010111000111111011;
		correct = 32'b00011001100010000000000101000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000101101011111100001001001;
		x2 = 32'b11101001111100000100111000110000;
		correct = 32'b01000000101100000100100000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000000101111101001000101101000;
		x2 = 32'b11011111110011010110010101111100;
		correct = 32'b11000000100011000000000101101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111011111001101011110011110111;
		x2 = 32'b00100010011000011100101111010100;
		correct = 32'b00100010011000001000100011010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101101101110011011111010101010;
		x2 = 32'b11101111100101001010101110101100;
		correct = 32'b10101101100100001010101010101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010000100011110100111011010001;
		x2 = 32'b01111110001000011010001001000011;
		correct = 32'b01010000000000010000001001000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001011111111101010001010100110;
		x2 = 32'b11100001010110110000011000010000;
		correct = 32'b00000001010110100000001000000000;
 #500; 
 			end  
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111001100010001001011001011;
		x2 = 32'b00000110001001111110110100101111;
		correct = 32'b00000110001000010000000000001011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011011010111000101001111111110;
		x2 = 32'b11100011000110011110100000100101;
		correct = 32'b00000011000110000100000000100100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100001111101011000100010000;
		x2 = 32'b01101001001100111000111110011101;
		correct = 32'b01101000001100101000000100010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100001110001011101101000010;
		x2 = 32'b01110100001110110000111001100111;
		correct = 32'b00010100001110000000101001000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101110001111001101100000101;
		x2 = 32'b01001111110111000001010001001011;
		correct = 32'b01000101110001000001000000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011111101010101110111010100001;
		x2 = 32'b00000001101000101110000011010101;
		correct = 32'b00000001101000101110000010000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001000010000010111111011100010;
		x2 = 32'b00110110101001011010100001010110;
		correct = 32'b00000000000000010010100001000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001001010001101000111010010101;
		x2 = 32'b01110010011001101100011100000010;
		correct = 32'b00000000010001101000011000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000000000100001001000111001100;
		x2 = 32'b11000011100001100011100011001110;
		correct = 32'b00000000000000000001000011001100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010010100100101100001000101111;
		x2 = 32'b10010011101011110101100100011111;
		correct = 32'b10010010100000100100000000001111;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001111000000110010111111101111;
		x2 = 32'b10100001111100101000010001010100;
		correct = 32'b00000001000000100000010001000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010101101100000011111001110101;
		x2 = 32'b01001001011110111001010000010100;
		correct = 32'b01000001001100000001010000010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001100000100010110100110111001;
		x2 = 32'b01110100101011110000001000101011;
		correct = 32'b00000100000000010000000000101001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110110010111001000110111011;
		x2 = 32'b10111101001110000000100011110110;
		correct = 32'b00111100000010000000000010110010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001001011010111011000001101100;
		x2 = 32'b10110010000000111111111010100010;
		correct = 32'b00000000000000111011000000100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001100110001111101001000011100;
		x2 = 32'b11100010101010001111011100100001;
		correct = 32'b01000000100000001101001000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101100010000000101001010101001;
		x2 = 32'b00111010101111010011011001101101;
		correct = 32'b00101000000000000001001000101001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011001010001111010000001110;
		x2 = 32'b00101101011101010100101010000000;
		correct = 32'b00000001001000000100000000000000;
 #500; 
 			end  
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111011001010111110011101101010;
		x2 = 32'b00100111010011001000101101001001;
		correct = 32'b00100011000010001000001101001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111010001010100111000101010010;
		x2 = 32'b11011100010111101011111111111000;
		correct = 32'b01011000000010100011000101010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111111100011111000101111011;
		x2 = 32'b10000000011001010010110011011100;
		correct = 32'b10000000011000010010000001011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010111001101001000101010011001;
		x2 = 32'b10100100010110010000000111101011;
		correct = 32'b10000100000100000000000010001001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110010000011101111100100010001;
		x2 = 32'b11001111110111011111110000110011;
		correct = 32'b11000010000011001111100000010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110001000100000011010001111100;
		x2 = 32'b11001110010111110101100101100011;
		correct = 32'b11000000000100000001000001100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010011100011110111111110011;
		x2 = 32'b10001001011010000110000111000111;
		correct = 32'b10001000011000000110000111000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011101110100000001101111111;
		x2 = 32'b11100010011111011100010001000010;
		correct = 32'b00100010001110000000000001000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011001111100110110010010001000;
		x2 = 32'b10011011000101000111011000100100;
		correct = 32'b10011001000100000110010000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110000010110110111011001011010;
		x2 = 32'b00011011000011011000011011001100;
		correct = 32'b00010000000010010000011001001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101010100110100001000110011111;
		x2 = 32'b11010001010011000100001010001000;
		correct = 32'b00000000000010000000000010001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000001100100111101110100110000;
		x2 = 32'b11101101001010101100100100011000;
		correct = 32'b00000001000000101100100100010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011011100110111100000110101;
		x2 = 32'b11000000011001000011101110100110;
		correct = 32'b01000000011000000011100000100100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010100001111011000111011000000;
		x2 = 32'b01010001111001000110011011011101;
		correct = 32'b00010000001001000000011011000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111100101111000100000101101;
		x2 = 32'b01011010101101010101000110011100;
		correct = 32'b00000010100101010000000000001100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100000111101101010100000010000;
		x2 = 32'b00111110000010001010010101001011;
		correct = 32'b00100000000000001010000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110011111101110110010111101100;
		x2 = 32'b01100011110101001001010010111011;
		correct = 32'b01100011110101000000010010101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011101111110101011100010111111;
		x2 = 32'b10101000100100000100101101100100;
		correct = 32'b10001000100100000000100000100100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000111001100000000111110011100;
		x2 = 32'b00111111010001000011010100001011;
		correct = 32'b00000111000000000000010100001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111111111001110010010000110010;
		x2 = 32'b10110111010111010111101100100110;
		correct = 32'b00110111010001010010000000100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000110100111010101100101110101;
		x2 = 32'b10010011011001011010001100001110;
		correct = 32'b10000010000001010000000100000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010001000011001000011101001010;
		x2 = 32'b10100000010100111101010001111011;
		correct = 32'b10000000000000001000010001001010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110000011110100101011010101;
		x2 = 32'b00101100010100111111001001101001;
		correct = 32'b00101100000000110100001001000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010110100100011111101101110100;
		x2 = 32'b01111110100010001110010110110000;
		correct = 32'b01010110100000001110000100110000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010010010000101101011100100011;
		x2 = 32'b01101000000111110101000101000011;
		correct = 32'b01000000000000100101000100000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001101100101111101001101110111;
		x2 = 32'b10101000101011010000100000110111;
		correct = 32'b10001000100001010000000000110111;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100111100111010010011001010101;
		x2 = 32'b10100111101110011110100101010110;
		correct = 32'b10100111100110010010000001010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011111100011111011111000110010;
		x2 = 32'b11011100011011011010011011001001;
		correct = 32'b00011100000011011010011000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011111000000011011010010010110;
		x2 = 32'b11111011111110001010100010111111;
		correct = 32'b10011011000000001010000010010110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000110000110000010000010001010;
		x2 = 32'b10100010111110111011011110001100;
		correct = 32'b10000010000110000010000010001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111011110101101010001011011100;
		x2 = 32'b00111001001000001101011101010010;
		correct = 32'b00111001000000001000001001010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111011011110110101100101010;
		x2 = 32'b00111110100110011000010000111000;
		correct = 32'b00110110000010010000000000101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101010001110110101111010011;
		x2 = 32'b00111010101101011101111101001010;
		correct = 32'b00100000000001010100101101000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011011001111110000010010001010;
		x2 = 32'b10000101111001010101000111110011;
		correct = 32'b10000001001001010000000010000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010000100011011101000011000000;
		x2 = 32'b00111000100111110111010101111100;
		correct = 32'b00010000100011010101000001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110110000010101110101001111;
		x2 = 32'b11011010101111101101100010001000;
		correct = 32'b00000010100000000101100000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110111010001100010000011001;
		x2 = 32'b11001111111100010010101001000000;
		correct = 32'b00000110111000000000000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011010000000001011000100000100;
		x2 = 32'b11111011001010110011100010111001;
		correct = 32'b11011010000000000011000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110010101010101011011110111101;
		x2 = 32'b01010111111011110000111101101010;
		correct = 32'b01010010101010100000011100101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110010000100110100111110000111;
		x2 = 32'b10100000000111010001000001010100;
		correct = 32'b10100000000100010000000000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100001111110010011101100010111;
		x2 = 32'b11110000011100110111101010010010;
		correct = 32'b01100000011100010011101000010010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001011001110101110100111011;
		x2 = 32'b00110111000110010110000110001111;
		correct = 32'b00110001000000010100000100001011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101110001010111101011000011011;
		x2 = 32'b10010000111101111000001100010111;
		correct = 32'b00000000001000111000001000010011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000011010000000001111100100;
		x2 = 32'b11100111010100101101100100101010;
		correct = 32'b10000000010000000000000100100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110110110011001110100001001001;
		x2 = 32'b01000001110001010010000110011100;
		correct = 32'b00000000110001000010000000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010100011100101001100111110101;
		x2 = 32'b10110010001010100111001100011111;
		correct = 32'b00010000001000100001000100010101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100011110110101110110101000111;
		x2 = 32'b10100101011011010010000110000100;
		correct = 32'b10100001010010000010000100000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101010101111011001110001101101;
		x2 = 32'b00000011000101101011011101000100;
		correct = 32'b00000010000101001001010001000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000110001011101010101110001001;
		x2 = 32'b10110011000101100010110011100100;
		correct = 32'b00000010000001100010100010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101010001000011000111100111;
		x2 = 32'b00100110100101110110010111101000;
		correct = 32'b00100100000001000010000111100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000111100000001000110101100;
		x2 = 32'b00011010010000001001100010101011;
		correct = 32'b00010000010000000001000010101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101000000001001000101110101010;
		x2 = 32'b11001010000110000010001111010100;
		correct = 32'b11001000000000000000001110000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111110011110010111000111111001;
		x2 = 32'b10011101100101100101000111100110;
		correct = 32'b10011100000100000101000111100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100000100100011100100101011;
		x2 = 32'b01111011100001111011110010010000;
		correct = 32'b01110000000000100011100000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100010100110001110100100110;
		x2 = 32'b10000100000011001110001111001110;
		correct = 32'b00000100000000000000000100000110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001101110000010001001011010;
		x2 = 32'b11010011000111100011011111010101;
		correct = 32'b00000001000110000010001001010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011010111111101010010110000010;
		x2 = 32'b01101011011110100110111101001000;
		correct = 32'b01001010011110100010010100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101000111110111101100000001010;
		x2 = 32'b01011100101110110000011000000001;
		correct = 32'b01001000101110110000000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111010100100011100000001000000;
		x2 = 32'b01001010000010101111010001100011;
		correct = 32'b01001010000000001100000001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011101101100010111000100111;
		x2 = 32'b10000010111011110010010010101010;
		correct = 32'b00000010101001100010010000100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011101101101110011000110011;
		x2 = 32'b11110100011101110010010101001001;
		correct = 32'b00100000001101100010010000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100100110000010001100100110110;
		x2 = 32'b01000000110100001111101111001000;
		correct = 32'b01000000110000000001100100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100101011001110111110000100110;
		x2 = 32'b00010011010100000110001001100000;
		correct = 32'b00000001010000000110000000100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111000001100111100110011101;
		x2 = 32'b11001101101111110011011101011001;
		correct = 32'b11000101000001100011000100011001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011011011100101011000101110010;
		x2 = 32'b10111010011100101100111010101011;
		correct = 32'b00011010011100101000000000100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101100010001010101101000011;
		x2 = 32'b00010011000110111110110101001100;
		correct = 32'b00000001000010001010100101000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010111010101010110000110011010;
		x2 = 32'b01011011010000110011110110001000;
		correct = 32'b00010011010000010010000110001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100111101100111011100101011111;
		x2 = 32'b10111111100011010111111100110001;
		correct = 32'b10100111100000010011100100010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011100110101101001000011110111;
		x2 = 32'b01111000110011010011101011011000;
		correct = 32'b00011000110001000001000011010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110100111010100001111100101111;
		x2 = 32'b00011101011001100011011010100110;
		correct = 32'b00010100011000100001011000100110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110000111000101100011011101100;
		x2 = 32'b00100000011111000011110010101111;
		correct = 32'b00100000011000000000010010101100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101011011101111100011011011;
		x2 = 32'b10101000011001001101000100110111;
		correct = 32'b00100000011001001101000000010011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000011001110111110110001110101;
		x2 = 32'b10110001000001001000011111000011;
		correct = 32'b00000001000000001000010001000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100110000101010110000110110001;
		x2 = 32'b01010000111100010111111111011100;
		correct = 32'b00000000000100010110000110010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001101011000110111100110101000;
		x2 = 32'b01101101010100101010000000000010;
		correct = 32'b00001101010000100010000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111011010001111101010101000;
		x2 = 32'b00101100011000110000101100101000;
		correct = 32'b00100100011000000000101000101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001100110001111101001000111011;
		x2 = 32'b00001111100100010100011100001001;
		correct = 32'b00001100100000010100001000001001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100000101011110000001011001111;
		x2 = 32'b00110011010001000001100011101011;
		correct = 32'b00100000000001000000000011001011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110000000011010010000010101101;
		x2 = 32'b10111101100110000110011011110011;
		correct = 32'b00110000000010000010000010100001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000001001110000101110101000;
		x2 = 32'b11011001000110010000011010100001;
		correct = 32'b10011000000000010000001010100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100011001000001001011001110;
		x2 = 32'b10100001001101110111001111010000;
		correct = 32'b10000000001001000001001011000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001110111011100101000010101010;
		x2 = 32'b00001111110001110011101001011110;
		correct = 32'b00001110110001100001000000001010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100001011111001111111010100;
		x2 = 32'b00100001110011010110001011000101;
		correct = 32'b00100000000011010000001011000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101001010101100111000111110111;
		x2 = 32'b00000000010011000101101101010001;
		correct = 32'b00000000010001000101000101010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000010100000100010101001010001;
		x2 = 32'b11110100110000101111011000111000;
		correct = 32'b00000000100000100010001000010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001110010000001000011110010101;
		x2 = 32'b10111101011100011110010100111111;
		correct = 32'b10001100010000001000010100010101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010110000111000100111110010000;
		x2 = 32'b11001100001110000010000010110001;
		correct = 32'b00000100000110000000000010010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011000001110111110111110000;
		x2 = 32'b00100011011011100000100010111100;
		correct = 32'b00000011000001100000100010110000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010010011111101111000111110010;
		x2 = 32'b10100100011111101011110001110000;
		correct = 32'b10000000011111101011000001110000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000001101011001111110101011001;
		x2 = 32'b00110111111001111100001011111010;
		correct = 32'b00000001101001001100000001011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101001001001000010100001011100;
		x2 = 32'b11000001001011111111010101111001;
		correct = 32'b01000001001001000010000001011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110001010101110001011000001;
		x2 = 32'b00110001001101000100110111000110;
		correct = 32'b00100000001000000100000011000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101111010111011011110011010;
		x2 = 32'b00111101110111100011011010001001;
		correct = 32'b00111101110010100011011010001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101011100000000111100110000000;
		x2 = 32'b00111110011001101001101010110001;
		correct = 32'b00101010000000000001100010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110000011010010011101111010001;
		x2 = 32'b01101101010000110011110000010001;
		correct = 32'b00100000010000010011100000010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100000010101100011110110100;
		x2 = 32'b01000001110001000000111101000001;
		correct = 32'b01000000000000000000011100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100010010011011000100111001111;
		x2 = 32'b00011100000000011110011001010110;
		correct = 32'b00000000000000011000000001000110;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100100000100111111111111111001;
		x2 = 32'b00110000111001000010110100000000;
		correct = 32'b00100000000000000010110100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000111100011001010011111010100;
		x2 = 32'b00110011001010100100011001000001;
		correct = 32'b00000011000010000000011001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000111101010010001010100100111;
		x2 = 32'b01101011001110011001001001000101;
		correct = 32'b01000011001010010001000000000101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010010100110111111010111100000;
		x2 = 32'b01100110011111111100100111101110;
		correct = 32'b01000010000110111100000111100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001110010111010110111100000;
		x2 = 32'b00010100111111100100101001011000;
		correct = 32'b00000000110010100000100001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110000011110110101000001101;
		x2 = 32'b01011100110100101101101011111000;
		correct = 32'b01011100000000100100101000001000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000101010100010001101010011;
		x2 = 32'b10111001111011110110001111100001;
		correct = 32'b10110000101010100010001101000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001000001011001010001011111011;
		x2 = 32'b11000110111000101110011101110111;
		correct = 32'b11000000001000001010001001110011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101001101000010000110011010;
		x2 = 32'b01110001100010011111101000110010;
		correct = 32'b01110001000000000010000000010010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110010100101110101110000001010;
		x2 = 32'b10011100010001011010110000110001;
		correct = 32'b00010000000001010000110000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100010111001001101111001011010;
		x2 = 32'b11000110100000010011010011110000;
		correct = 32'b01000010100000000001010001010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011110101110000011101011011001;
		x2 = 32'b11110000011010100111001110111110;
		correct = 32'b01010000001010000011001010011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101001000000011110001010000110;
		x2 = 32'b10001100100100000110101110010100;
		correct = 32'b10001000000000000110001010000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101011101011101111000011101000;
		x2 = 32'b00010101011001111101100011010100;
		correct = 32'b00000001001001101101000011000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100100100111001000111110100010;
		x2 = 32'b10111001001101011111101110111000;
		correct = 32'b00100000000101001000101110100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101011001000010101001011001010;
		x2 = 32'b01000101110101011000001110100010;
		correct = 32'b00000001000000010000001010000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101100111001001110100111101111;
		x2 = 32'b00000011101001011001101101110010;
		correct = 32'b00000000101001001000100101100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100011000010011110011010010001;
		x2 = 32'b10010101010010101110111011100010;
		correct = 32'b10000001000010001110011010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111001010111011101101101000111;
		x2 = 32'b00001100000000100000011010111100;
		correct = 32'b00001000000000000000001000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111000000111110111101010111011;
		x2 = 32'b10000111010110111010111001011100;
		correct = 32'b00000000000110110010101000011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100010001010111111111100010010;
		x2 = 32'b01011100110100001110111010010000;
		correct = 32'b01000000000000001110111000010000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100001010100100010001101110101;
		x2 = 32'b00000010011110000001011110011100;
		correct = 32'b00000000010100000000001100010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011000011010001000111000011000;
		x2 = 32'b00101011000101101011010001111111;
		correct = 32'b00001000000000001000010000011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001111010110100001000011001100;
		x2 = 32'b01011101010010101101001110101110;
		correct = 32'b01001101010010100001000010001100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011000011001001100010111101010;
		x2 = 32'b00110011010110100111010011000100;
		correct = 32'b00010000010000000100010011000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100100010011010011000011101100;
		x2 = 32'b11001100111100100011001111000111;
		correct = 32'b00000100010000000011000011000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111100100011001110100011101010;
		x2 = 32'b00100101000111111101000110010111;
		correct = 32'b00100100000011001100000010000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011111111100011001010011101;
		x2 = 32'b11000011101111110001101101110011;
		correct = 32'b10000011101111100001001000010001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111110101100000011011010001001;
		x2 = 32'b00001101101011010110110110100101;
		correct = 32'b00001100101000000010010010000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001100111010001110100101100;
		x2 = 32'b00011111010000110001010110010010;
		correct = 32'b00000001000000010001010100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101001000010011011001101111111;
		x2 = 32'b11000000111111000000110111010111;
		correct = 32'b11000000000010000000000101010111;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001001011010101100000110011000;
		x2 = 32'b11100000101010100001100010011110;
		correct = 32'b11000000001010100000000010011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100100011100000110100011011001;
		x2 = 32'b10001011010100110001100001011000;
		correct = 32'b10000000010100000000100001011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010110101001001010001001100010;
		x2 = 32'b10010101100110100010011001111110;
		correct = 32'b10010100100000000010001001100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000011110110011110100001000010;
		x2 = 32'b10011011111110111010101100100100;
		correct = 32'b00000011110110011010100000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110111001100110010000011010000;
		x2 = 32'b11010001001011100101100011101100;
		correct = 32'b10010001001000100000000011000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100110101001100001010111001011;
		x2 = 32'b00000011101110100101111101000111;
		correct = 32'b00000010101000100001010101000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101011101001010101111011000;
		x2 = 32'b00110011000110101110011001100010;
		correct = 32'b00100001000100001010001001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000010101010100101110101110111;
		x2 = 32'b10100111101000000111101010111100;
		correct = 32'b00000010101000000101100000110100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001100011101011011111101110011;
		x2 = 32'b11101010000101111010010011000010;
		correct = 32'b00001000000101011010010001000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111101111001010101010001000100;
		x2 = 32'b00010001000001110001010111000011;
		correct = 32'b00010001000001010001010001000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100111001011000011100000001111;
		x2 = 32'b11010101101110111010011001100100;
		correct = 32'b01000101001010000010000000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110101001011001101001101000100;
		x2 = 32'b10101110100001101100100110110111;
		correct = 32'b10100100000001001100000100000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010011011111010001011000111001;
		x2 = 32'b10101001000101011011101011000001;
		correct = 32'b10000001000101010001001000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111011100110110011000010101;
		x2 = 32'b10001110001010010101001010100011;
		correct = 32'b00000110001000010100001000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011111101000110000110110111011;
		x2 = 32'b00100101101010111000001111101011;
		correct = 32'b00000101101000110000000110101011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011111011110001110001000001100;
		x2 = 32'b01100110000000011000001000000010;
		correct = 32'b00000110000000001000001000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101010010010000111110110111000;
		x2 = 32'b01001000100110110011101101101001;
		correct = 32'b00001000000010000011100100101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101101011101100011111000101;
		x2 = 32'b00100001011101011011110100000111;
		correct = 32'b00100001001001001000010100000101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010000110001101010000010011000;
		x2 = 32'b11011011100111001111100110000111;
		correct = 32'b11010000100001001010000010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111001011100100110010000000;
		x2 = 32'b11100010000100010110001001000000;
		correct = 32'b00100010000000000100000000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011101100010101111001010010;
		x2 = 32'b11101001001010000000110110000111;
		correct = 32'b01001001001000000000110000000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111111101010111001101110101;
		x2 = 32'b01001011111111000111100011000001;
		correct = 32'b00000011111101000111000001000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010111000110011110010101110;
		x2 = 32'b11110001000011001011111111010000;
		correct = 32'b01000000000000000011110010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010100000111000010011011011011;
		x2 = 32'b01111101010101100010111000100111;
		correct = 32'b01010100000101000010011000000011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111100011000110000111011010101;
		x2 = 32'b10011100110100001110010101000011;
		correct = 32'b00011100010000000000010001000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100111000000000101110110110010;
		x2 = 32'b11011001011010010110101101111101;
		correct = 32'b11000001000000000100100100110000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100001000100011101011010011100;
		x2 = 32'b00001100001110100000001110111000;
		correct = 32'b00000000000100000000001010011000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101000010011010011011011000101;
		x2 = 32'b00111110100010010001101110001100;
		correct = 32'b00101000000010010001001010000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011111111101111000100110000011;
		x2 = 32'b01111011110000111010010100010110;
		correct = 32'b01011011110000111000000100000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100110001111000001110111001110;
		x2 = 32'b01010101101011101001000110010000;
		correct = 32'b01000100001011000001000110000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111010000101000110100110000;
		x2 = 32'b11100001001101111101011001001011;
		correct = 32'b11000001000000101000010000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011011011101101001100000000111;
		x2 = 32'b01000001101001000000110000001000;
		correct = 32'b01000001001001000000100000000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111111000110000011110110111111;
		x2 = 32'b10001001011001001000000010000000;
		correct = 32'b00001001000000000000000010000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100000110100011110010110010110;
		x2 = 32'b10100111111101010000101110001011;
		correct = 32'b10100000110100010000000110000010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001000111000011000001101100001;
		x2 = 32'b01101111101111110111000101110010;
		correct = 32'b00001000101000010000000101100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000100101101000001011100111010;
		x2 = 32'b00101000000000110110010110101100;
		correct = 32'b00000000000000000000010100101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100001111111000010100011101;
		x2 = 32'b00010011010110111100100110010100;
		correct = 32'b00010000000110111000000100010100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111101101100010011010101110;
		x2 = 32'b11001111111111110111100111110001;
		correct = 32'b10001111101101100010000010100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111010000010011111001100101011;
		x2 = 32'b11000110001011111110011110100110;
		correct = 32'b11000010000010011110001100100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001011001101110110011011110;
		x2 = 32'b01011111111000001111110001100100;
		correct = 32'b00000001011000001110110001000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110011101101101100010001110101;
		x2 = 32'b00011000100000111100000101111100;
		correct = 32'b00010000100000101100000001110100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101111000100100111001111101110;
		x2 = 32'b01111111111101111100011101110001;
		correct = 32'b00101111000100100100001101100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110111100010010101001100010011;
		x2 = 32'b11001111011100100000011101100101;
		correct = 32'b11000111000000000000001100000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001101111010100101100101001111;
		x2 = 32'b11011011011101101111010011001011;
		correct = 32'b00001001011000100101000001001011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101101001110010110111110100100;
		x2 = 32'b11000000100001111010010001000100;
		correct = 32'b10000000000000010010010000000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101011011100001011110001100101;
		x2 = 32'b00000101010000010100111101111110;
		correct = 32'b00000001010000000000110001100100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111011110000000011001011111;
		x2 = 32'b10001100011110001000110110111111;
		correct = 32'b10001100011110000000010000011111;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011100001011100101001001000101;
		x2 = 32'b01010001011000001111111101011011;
		correct = 32'b01010000001000000101001001000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110100111010011001100001100;
		x2 = 32'b01111101110111110101001111101101;
		correct = 32'b00000100100111010001001100001100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100100011011110000110000001101;
		x2 = 32'b00011101010100011011010000101001;
		correct = 32'b00000100010000010000010000001001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011100000111100110101101001110;
		x2 = 32'b10111111100001110011001110010000;
		correct = 32'b00011100000001100010001100000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001000110110111110011001011011;
		x2 = 32'b10000111001111100000110101001111;
		correct = 32'b00000000000110100000010001001011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011001001001011101111001110110;
		x2 = 32'b01101010101111011001100001100011;
		correct = 32'b00001000001001011001100001100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010000110100000001111010111010;
		x2 = 32'b00011000100010110011000111100010;
		correct = 32'b00010000100000000001000010100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011101001000011111011111000001;
		x2 = 32'b10111001110001100001011111100110;
		correct = 32'b00011001000000000001011111000000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001110100001000011100000010011;
		x2 = 32'b10001001101000000110000010001001;
		correct = 32'b10001000100000000010000000000001;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000101011000110001100011100100;
		x2 = 32'b10100100010000001101101101001111;
		correct = 32'b00000100010000000001100001000100;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010011010101011111001011100010;
		x2 = 32'b10001101000111110111110010111001;
		correct = 32'b00000001000101010111000010100000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001101111001111011110010100010;
		x2 = 32'b10000110101000010001010001110111;
		correct = 32'b00000100101000010001010000100010;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101001010000101001110111011;
		x2 = 32'b01010001111001111100101011110011;
		correct = 32'b00010001001000000100001010110011;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011101110011001011011000010111;
		x2 = 32'b01101111010011100110110000000101;
		correct = 32'b00001101010011000010010000000101;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011100100010011011100011111110;
		x2 = 32'b10100011101000111000111111111001;
		correct = 32'b10000000100000011000100011111000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101110100100000101011111111100;
		x2 = 32'b11000001111011111000000101101001;
		correct = 32'b01000000100000000000000101101000;
 #500; 
 			end 
 begin
			$display ("x1      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("x2      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("x3 : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end
end 
endmodule