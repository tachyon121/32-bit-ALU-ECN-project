`timescale 1 ns/1 ps
    `include "alu.v"


    module mul_tb ();
        reg clock;
        reg [31:0] x1, x2;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] x3;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .x1(x1),
                .x2(x2),
                .OpCode(op),
                .x3(x3)
            );
        /* create x1 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, x1, x2, op, x3);
            clock = 0;

    op = 3'b011;

		/* Display the operation */
		$display ("Opcode: 011, Operation: MUL");
		/* Test Cases!*/
		x1 = 32'b00001001111010001000001111111101;
		x2 = 32'b01101111100001111011001011000110;
		correct = 32'b00111001111101100111111111110100;
		#400; //5.597609e-33 * 8.39932e+28 = 0.0004701611
					
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011110011010110001111101001100;
		x2 = 32'b11000100100010001000010100100000;
		correct = 32'b01100011011110101100010111001010;
		#400; //-4.235586e+18 * -1092.1602 = 4.6259382e+21
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110011010000110000001010100;
		x2 = 32'b11010010111000010100010010100110;
		correct = 32'b10011001110011000111101011111010;
		#400; //4.370512e-35 * -483759700000.0 = -2.1142775e-23
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111111111011110010111100110000;
		x2 = 32'b01110000000000100101001100001010;
		correct = 32'b11111111111011110010111100110000;
		#400; //nan * 1.6133376e+29 = nan
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101101010000011100101111011100;
		x2 = 32'b10111100000001010001010001111001;
		correct = 32'b10101001110010010111110011010010;
		#400; //1.1016046e-11 * -0.008122557 = -8.947846e-14
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110000010111101111001110010100;
		x2 = 32'b11001101111111100011101001101011;
		correct = 32'b11111110110111010110100010001101;
		#400; //2.7600056e+29 * -533155170.0 = -1.4715112e+38
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111110111000111100010011000010;
		x2 = 32'b11100111001110010001001110111111;
		correct = 32'b01100110101001001010101011000010;
		#400; //-0.44486052 * -8.7400205e+23 = 3.88809e+23
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101010010011010010111111010101;
		x2 = 32'b11110100101100111011011111011000;
		correct = 32'b01011111100100000000101111001100;
		#400; //-1.8224253e-13 * -1.139099e+32 = 2.0759228e+19
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010101111001010110111100010100;
		x2 = 32'b11010011101111100101011111001110;
		correct = 32'b10101010001010101001011100100010;
		#400; //9.2667614e-26 * -1635033800000.0 = -1.5151468e-13
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000110111100111101000111111001;
		x2 = 32'b11110011011111100011011110011101;
		correct = 32'b01111010111100100001111101001101;
		#400; //-31208.986 * -2.0141165e+31 = 6.2858535e+35
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001010000101111011100011111011;
		x2 = 32'b00111011110101001111010110111110;
		correct = 32'b10000110011111000110110110101001;
		#400; //-7.3051765e-33 * 0.0064990213 = -4.7476498e-35
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101001001011000101001011111000;
		x2 = 32'b00010010001010001011111010100011;
		correct = 32'b10111011111000110010110110001100;
		#400; //-1.3020441e+25 * 5.324643e-28 = -0.00693292
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100101101001001111110000111010;
		x2 = 32'b01000100011110111101111011100000;
		correct = 32'b01101010101000100101001011110000;
		#400; //9.739011e+22 * 1007.4824 = 9.811882e+25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101000011001000101100111101010;
		x2 = 32'b11000000101101101001010100111001;
		correct = 32'b00101001101000101101110100001000;
		#400; //-1.26760395e-14 * -5.7057157 = 7.232588e-14
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010111011001100010101101000000;
		x2 = 32'b11100100100001101110000001111100;
		correct = 32'b10111100011100101000100011110010;
		#400; //7.4371597e-25 * -1.9904316e+22 = -0.014803158
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111100110010001100110000110010;
		x2 = 32'b10100011000010100011110000110000;
		correct = 32'b11100000010110001101101010010001;
		#400; //8.3408076e+36 * -7.49374e-18 = -6.2503845e+19
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010111010111011100010001100110;
		x2 = 32'b11011000011010110000110011111010;
		correct = 32'b11110000010010111001111010000111;
		#400; //243835600000000.0 * -1033763870000000.0 = -2.5206842e+29
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000101011011111010001110111;
		x2 = 32'b01001101001011100101000011010001;
		correct = 32'b10100110011011001110011000100111;
		#400; //-4.49663e-24 * 182783250.0 = -8.2190863e-16
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100101011101110011011001101110;
		x2 = 32'b01000110010011111000011110101111;
		correct = 32'b01101100010010000110100000001010;
		#400; //7.2964286e+22 * 13281.921 = 9.691059e+26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010001011010010010001011000000;
		x2 = 32'b01000000000100011000011110111110;
		correct = 32'b00010010000001001000100001001101;
		#400; //1.8391167e-28 * 2.27391 = 4.181986e-28
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111001110111000110011100010000;
		x2 = 32'b01000010011101111010001110111110;
		correct = 32'b10111100110101010011010001101010;
		#400; //-0.00042038457 * 61.909904 = -0.02602597
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110000100010011111011000111101;
		x2 = 32'b00101101011100010100110000001001;
		correct = 32'b00011110100000100000100111001001;
		#400; //1.0038047e-09 * 1.3716147e-11 = 1.3768332e-20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011010111010111000000100011011;
		x2 = 32'b00110101001110000001000101100001;
		correct = 32'b00010000101010010101010011001000;
		#400; //9.74023e-23 * 6.857063e-07 = 6.678937e-29
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000100011100011100111000111110;
		x2 = 32'b11101000111100000011101001100110;
		correct = 32'b00101101111000101110100010000011;
		#400; //-2.8424116e-36 * -9.075562e+24 = 2.5796481e-11
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110000010111001111100100001010;
		x2 = 32'b10100101010000110000110110001100;
		correct = 32'b00010110001010000101110101100100;
		#400; //-8.038944e-10 * -1.6918144e-16 = 1.3600401e-25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000111001010010100101011010;
		x2 = 32'b10000101000101111000010001110101;
		correct = 32'b10010110100001111010000111110110;
		#400; //30757540000.0 * -7.1243144e-36 = -2.1912638e-25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101100101011010011010100011001;
		x2 = 32'b00101000100111011010010000000011;
		correct = 32'b10010101110101010101000100010001;
		#400; //-4.9228508e-12 * 1.750163e-14 = -8.6157915e-26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101110011001010110100101110;
		x2 = 32'b00111010110000011111101100111001;
		correct = 32'b00000001000110110001011101101011;
		#400; //1.9247684e-35 * 0.0014799602 = 2.8485805e-38
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011011101001101001110010100010;
		x2 = 32'b01001101111010001010111111100101;
		correct = 32'b01101010000101110111000001101101;
		#400; //9.379413e+16 * 487980200.0 = 4.576968e+25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000110001011000000111000111101;
		x2 = 32'b01100000100011010001010110000011;
		correct = 32'b11100111001111011010010010011010;
		#400; //-11011.56 * 8.132941e+19 = -8.955636e+23
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110010000000001110100010011011;
		x2 = 32'b10100011100101110001101111110100;
		correct = 32'b11010110000110000010111010001110;
		#400; //2.5532982e+30 * -1.6383291e-17 = -41831430000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000110011010100101000111100011;
		x2 = 32'b00101111110000010101101100110101;
		correct = 32'b10110110101100001111101100111000;
		#400; //-14996.472 * 3.5171302e-10 = -5.2744545e-06
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011011100111110101011000110001;
		x2 = 32'b01001010111001111100000011011011;
		correct = 32'b10100111000100000011111011001111;
		#400; //-2.6360043e-22 * 7594093.5 = -2.0018063e-15
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100111111011000111100010001111;
		x2 = 32'b11110110011011001100111101101011;
		correct = 32'b01011110110110101011111010111100;
		#400; //-6.563387e-15 * -1.2007705e+33 = 7.881121e+18
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010011001000110111010111000101;
		x2 = 32'b01100011000010100001100001101010;
		correct = 32'b11110110101100000101101000100110;
		#400; //-702055500000.0 * 2.54741e+21 = -1.7884232e+33
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100100100111011000101101100;
		x2 = 32'b01111101000000110101000010000101;
		correct = 32'b11010010000101111000010001111101;
		#400; //-1.4913187e-26 * 1.0909184e+37 = -162690710000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100110000110111111011100111000;
		x2 = 32'b11110100110111001111101010101001;
		correct = 32'b01011011100001101010000100101011;
		#400; //-5.411147e-16 * -1.4006217e+32 = 7.578971e+16
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100001010001011011111111111111;
		x2 = 32'b00100000000000110101001000101101;
		correct = 32'b00000001110010101110000101110011;
		#400; //6.70003e-19 * 1.1123321e-19 = 7.4526585e-38
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100000001010101010100000111;
		x2 = 32'b10111010110000010111111111010001;
		correct = 32'b00110111010010011000111101011001;
		#400; //-0.008137948 * -0.0014762824 = 1.2013909e-05
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100110000001111111111111110100;
		x2 = 32'b11000101011111101011110100010111;
		correct = 32'b01101100000001110101010001101000;
		#400; //-1.6056024e+23 * -4075.818 = 6.544143e+26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001000001110110010111111000100;
		x2 = 32'b10101100001010111001101100110010;
		correct = 32'b10110100111110101111010011000101;
		#400; //191679.06 * -2.4386712e-12 = -4.6744222e-07
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111100011011011001111010001;
		x2 = 32'b11000110101010110001001100100100;
		correct = 32'b10101110101111010110001101101010;
		#400; //3.933032e-15 * -21897.57 = -8.6123844e-11
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001010010000110111011001110100;
		x2 = 32'b01011000110010010011010011101110;
		correct = 32'b11100011100110011010000001101011;
		#400; //-3202461.0 * 1769833300000000.0 = -5.6678224e+21
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110101000010000100011000110110;
		x2 = 32'b10111101100110011000111100010100;
		correct = 32'b11110011001000110111110001000000;
		#400; //1.7274815e+32 * -0.07497993 = -1.2952644e+31
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001001111100000011101001111011;
		x2 = 32'b00111101110101010001111000111110;
		correct = 32'b00001000010001111111110100001001;
		#400; //5.7832893e-33 * 0.10406159 = 6.0181826e-34
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111110110101010111100110011001;
		x2 = 32'b00100000000100001001110101110011;
		correct = 32'b01011111011100010010111101100011;
		#400; //1.4187847e+38 * 1.224937e-19 = 1.7379218e+19
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101111000110111100101011100101;
		x2 = 32'b01001100010110111001010001011111;
		correct = 32'b01111100000001011010000011011101;
		#400; //4.821546e+28 * 57561468.0 = 2.7753527e+36
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110110001011101010110000100011;
		x2 = 32'b00000100111101110110100111010001;
		correct = 32'b10111011101010001101000001001001;
		#400; //-8.856943e+32 * 5.8166598e-36 = -0.0051517827
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001100010101011110111011111010;
		x2 = 32'b01111101010000000000001011100011;
		correct = 32'b01001010001000000111010110100101;
		#400; //1.6480838e-31 * 1.5951673e+37 = 2628969.2
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001010110100111111101110000111;
		x2 = 32'b11111010111111110011100000111110;
		correct = 32'b01000110010100110101011000011110;
		#400; //-2.0413175e-32 * -6.625882e+35 = 13525.529
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011011000010110111110001101001;
		x2 = 32'b11111010111001011000010010101001;
		correct = 32'b11010110011110100001110100100100;
		#400; //1.153801e-22 * -5.9586332e+35 = -68750766000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010001011110011001110001011100;
		x2 = 32'b11101110101000000011111100000000;
		correct = 32'b01000000100111000011111100100111;
		#400; //-1.9690818e-28 * -2.4796882e+28 = 4.882709
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011111000000001011101101101110;
		x2 = 32'b10000001100000100010110111101011;
		correct = 32'b10100001000000101110110010001010;
		#400; //9.276129e+18 * -4.7820347e-38 = -4.435877e-19
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101010100010001000100001100001;
		x2 = 32'b10110001111010110111000101010110;
		correct = 32'b11011100111110110010001101000110;
		#400; //8.252897e+25 * -6.852285e-09 = -5.6551202e+17
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000101110101000101100110111001;
		x2 = 32'b01001110011111100011001011111101;
		correct = 32'b11010100110100101101101101010001;
		#400; //-6795.2153 * 1066188600.0 = -7244981000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001101110001000111100111011111;
		x2 = 32'b01000000101010101010100111111011;
		correct = 32'b11001111000000101111101101100011;
		#400; //-412040160.0 * 5.3332496 = -2197513000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000111111010000010000011001100;
		x2 = 32'b01010010011011010101111001000000;
		correct = 32'b10011010110101110011101111010011;
		#400; //-3.4926757e-34 * 254872130000.0 = -8.901857e-23
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001100100101101110111100101;
		x2 = 32'b01110010011100111101001010010100;
		correct = 32'b01011100100010111110000101101111;
		#400; //6.522195e-14 * 4.8294036e+30 = 3.149831e+17
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110011100010000001110101110101;
		x2 = 32'b11000001000001001010001101011101;
		correct = 32'b01110101000011010000110000011001;
		#400; //-2.1568293e+31 * -8.289884 = 1.7879864e+32
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001011000000101001101011101010;
		x2 = 32'b01101000100010010001000111010000;
		correct = 32'b11110100000010111101101111111011;
		#400; //-8559338.0 * 5.1783423e+24 = -4.432318e+31
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001011100011011010111001001;
		x2 = 32'b01101010110010010011010011000001;
		correct = 32'b01010100101111011111100110001010;
		#400; //5.3670423e-14 * 1.2162161e+26 = 6527483000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010110000010001111001101010110;
		x2 = 32'b01100101011110101010010000100010;
		correct = 32'b10111100000001100001010101110000;
		#400; //-1.1062776e-25 * 7.397621e+22 = -0.008183822
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110000011001010000100111010100;
		x2 = 32'b00111000100100011011101000000010;
		correct = 32'b11101001100000100110000011111100;
		#400; //-2.835358e+29 * 6.9487854e-05 = -1.9702294e+25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110101010001010001100111111;
		x2 = 32'b11010110111001101010100001110010;
		correct = 32'b10111110000101111111000110100001;
		#400; //1.170159e-15 * -126805570000000.0 = -0.14838268
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110111000001110101010000110;
		x2 = 32'b01111001110110000100100001100110;
		correct = 32'b01000001001111100000010101111101;
		#400; //8.4604036e-35 * 1.4037557e+35 = 11.87634
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100011011100001111110001101011;
		x2 = 32'b11101110111010110101010101111100;
		correct = 32'b01010010110111011000100000101111;
		#400; //-1.3063878e-17 * -3.641616e+28 = 475736280000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111101000101110001100011101111;
		x2 = 32'b01111011110110110110000000100000;
		correct = 32'b11111001100000010111101100010001;
		#400; //-0.036889013 * 2.2781253e+36 = -8.40378e+34
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100001100111010000111110111;
		x2 = 32'b10011000101101110110110011111010;
		correct = 32'b00010101100000001011010100111111;
		#400; //-0.010963908 * -4.741443e-24 = 5.1984744e-26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100010011110001001010101011110;
		x2 = 32'b01100101011000001011110001101010;
		correct = 32'b01001000010110100011100110100111;
		#400; //3.3689342e-18 * 6.6330357e+22 = 223462.61
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100010001101111110000100111001;
		x2 = 32'b00011000001001000010011010010111;
		correct = 32'b00111010111010111101000000000001;
		#400; //8.479958e+20 * 2.1215986e-24 = 0.0017991067
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111101111010001010011011010011;
		x2 = 32'b10101101000111101111110100101101;
		correct = 32'b11101011100100000111110100001100;
		#400; //3.8655887e+37 * -9.0374765e-12 = -3.4935167e+26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110010100001101000011000110000;
		x2 = 32'b10010111010011110111001001000101;
		correct = 32'b11001010010110100000010100011010;
		#400; //5.3290514e+30 * -6.7029536e-25 = -3572038.5
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100000010111010100000001100111;
		x2 = 32'b10100110110100001000000001110110;
		correct = 32'b11000111101101000011001101011010;
		#400; //6.3771424e+19 * -1.4467719e-15 = -92262.7
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011101110110010001010110110;
		x2 = 32'b11010001010111010101111100111011;
		correct = 32'b10110101101000011101001010010100;
		#400; //2.0289281e-17 * -59424092000.0 = -1.2056721e-06
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101011110001101100111011001011;
		x2 = 32'b00100110011000110110100101110100;
		correct = 32'b11010010101100001001101101000011;
		#400; //-4.8068773e+26 * 7.889936e-16 = -379259550000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001101010010100001110111100011;
		x2 = 32'b11101010111110101001000100101000;
		correct = 32'b01111000110001011101001111001010;
		#400; //-211934770.0 * -1.5145847e+26 = 3.2099315e+34
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001101010111100000100001111;
		x2 = 32'b00100101111011001000100001100111;
		correct = 32'b01100000000111101011000101111101;
		#400; //1.1147481e+35 * 4.1031904e-16 = 4.5740233e+19
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101010100100110101111101100011;
		x2 = 32'b00010010011110011010110010101111;
		correct = 32'b00111101100011111011101100110000;
		#400; //8.908127e+25 * 7.8783395e-28 = 0.07018125
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000111101011101011110101110101;
		x2 = 32'b00010101001000110110010001100001;
		correct = 32'b00011101010111110000111001001011;
		#400; //89466.914 * 3.2996773e-26 = 2.9521194e-21
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100011011000101010110010010001;
		x2 = 32'b11010110100111000000101001001011;
		correct = 32'b01111010100010100010101001000110;
		#400; //-4.181399e+21 * -85784010000000.0 = 3.586972e+35
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010001001100001111110000001100;
		x2 = 32'b11110111100101011001010100001101;
		correct = 32'b01001001010011101101001101111101;
		#400; //-1.396162e-28 * -6.067776e+33 = 847159.8
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101110100011001010001111111;
		x2 = 32'b00111100011001111100110101000001;
		correct = 32'b00000010101111011100010100001000;
		#400; //1.9708814e-35 * 0.014148057 = 2.7884144e-37
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111001011111010100011000000100;
		x2 = 32'b10011011010000111010100010101010;
		correct = 32'b01010101010000011001001100110011;
		#400; //-8.219195e+34 * -1.618452e-22 = 13302372000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010011000010000010100011100;
		x2 = 32'b10000110100110000101101110100000;
		correct = 32'b10001001100001011110101110010010;
		#400; //56.25499 * -5.7310676e-35 = -3.2240115e-33
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100100001011100110111111110;
		x2 = 32'b01001000010000100010110100011110;
		correct = 32'b01111101010010101111101101011111;
		#400; //8.480878e+31 * 198836.47 = 1.6863078e+37
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100000000101010101010100001010;
		x2 = 32'b11000111010000110110111110100100;
		correct = 32'b10100111111001000000000111001100;
		#400; //1.2648928e-19 * -50031.64 = -6.328466e-15
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111001101111011111101110111011;
		x2 = 32'b00001110111101001011110100011000;
		correct = 32'b00001001001101011010000001000011;
		#400; //0.00036236443 * 6.0332735e-30 = 2.1862437e-33
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000010011100100001011000010101;
		x2 = 32'b01110101110110110000110010000111;
		correct = 32'b11111000110011110010010010111101;
		#400; //-60.521564 * 5.5535503e+32 = -3.3610956e+34
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101101100100000010111110110011;
		x2 = 32'b00100111001111111010111101111011;
		correct = 32'b00010101010101111110110011011001;
		#400; //1.6392087e-11 * 2.6601703e-15 = 4.3605744e-26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111111110111011101100001011010;
		x2 = 32'b10101010100111001000000101011110;
		correct = 32'b00101011000001111001111111110010;
		#400; //-1.733165 * -2.7800933e-13 = 4.8183603e-13
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010110101100000111101101010000;
		x2 = 32'b00010101111000101110001001101111;
		correct = 32'b00101101000111000110100011110110;
		#400; //97021835000000.0 * 9.163792e-26 = 8.890879e-12
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000110011001010001010010001001;
		x2 = 32'b00111011011100100000110001101111;
		correct = 32'b11000010010110001001100010001010;
		#400; //-14661.134 * 0.003693368 = -54.148964
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100100010101001010101001001101;
		x2 = 32'b10101001100000000000001110110101;
		correct = 32'b00001110010101001011000001110110;
		#400; //-4.6114422e-17 * -5.684985e-14 = 2.621598e-30
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110011010001100010100111100001;
		x2 = 32'b00111111010101101011000110110111;
		correct = 32'b10110011001001100011000010010011;
		#400; //-4.6138556e-08 * 0.8386492 = -3.8694065e-08
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011001100011010010100100100010;
		x2 = 32'b00110101111111100001011011111010;
		correct = 32'b01010000000011000001101101111011;
		#400; //4966649700000000.0 * 1.8931162e-06 = 9402445000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011110100000101111010101110001;
		x2 = 32'b01111010001001110010100101111000;
		correct = 32'b01011001001010110000011010100111;
		#400; //1.3865798e-20 * 2.1698867e+35 = 3008721000000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111000111000010110101010111;
		x2 = 32'b00010001010010010100001010000011;
		correct = 32'b10101000111101011001000001011010;
		#400; //-171718550000000.0 * 1.58766e-28 = -2.7263067e-14
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000000010101001110010000011;
		x2 = 32'b00001100000001110100011101011101;
		correct = 32'b00011100100100100111111001011010;
		#400; //9302052000.0 * 1.0421497e-31 = 9.694131e-22
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111011100001011001110010101101;
		x2 = 32'b10111000000110000010010001100001;
		correct = 32'b00110100000111101101000000000111;
		#400; //-0.004077515 * -3.6273505e-05 = 1.4790577e-07
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100000010010010111100001111;
		x2 = 32'b10100010110010100101110101110100;
		correct = 32'b00110111010110001110001001101100;
		#400; //-2356800000000.0 * -5.4851157e-18 = 1.2927321e-05
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001011010111001011100111101110;
		x2 = 32'b01100010101000110011011010000001;
		correct = 32'b10101110100011001011100101100001;
		#400; //-4.2510337e-32 * 1.5053734e+21 = -6.399393e-11
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111100011110010101001111110;
		x2 = 32'b01111101011101011100001010111000;
		correct = 32'b01110101100010010111000010010000;
		#400; //1.7066715e-05 * 2.0416994e+37 = 3.4845103e+32
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000101101100001001010011110100;
		x2 = 32'b01110110110101010011110101101010;
		correct = 32'b00111101000100110001011001001100;
		#400; //1.6605677e-35 * 2.1625095e+33 = 0.035909936
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100011001100011101101011101110;
		x2 = 32'b00010001111001110010110000010111;
		correct = 32'b00110101101000001001101100101110;
		#400; //3.2808492e+21 * 3.6472546e-28 = 1.1966092e-06
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100110100011110000100110101000;
		x2 = 32'b01001011010100101000011010011110;
		correct = 32'b00110010011010110100001001000110;
		#400; //9.925236e-16 * 13797022.0 = 1.3693869e-08
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011011101100010010100010110001;
		x2 = 32'b01010101010110100011111111000100;
		correct = 32'b11110001100101110000100011000111;
		#400; //-9.973162e+16 * 14997963000000.0 = -1.4957711e+30
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011001110111110110111110100100;
		x2 = 32'b10100011011101110001111101100010;
		correct = 32'b00111101110101111011000000011011;
		#400; //-7861459000000000.0 * -1.3396542e-17 = 0.10531636
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100100100110010000100011010000;
		x2 = 32'b11010100101111100011100111011101;
		correct = 32'b01111001111000110110111001000011;
		#400; //-2.2583895e+22 * -6536116600000.0 = 1.4761097e+35
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011000110101110010001011000111;
		x2 = 32'b00110100010000011101000101110000;
		correct = 32'b00001101101000101110000100111010;
		#400; //5.5611314e-24 * 1.8050719e-07 = 1.0038242e-30
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000111000011110010101110011;
		x2 = 32'b01000000110000100000110110101000;
		correct = 32'b01010010001010110011101111101110;
		#400; //30319286000.0 * 6.064167 = 183861220000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101000111000001000111011010;
		x2 = 32'b11000011001011001001111011000000;
		correct = 32'b00101000110100100111100110001101;
		#400; //-1.3536891e-16 * -172.62012 = 2.3367398e-14
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000110111010100011101000010011;
		x2 = 32'b11011110001010000110011001011011;
		correct = 32'b10100101100110100001001111000011;
		#400; //8.810635e-35 * -3.0336216e+18 = -2.6728133e-16
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000010001011010001011010100110;
		x2 = 32'b10111111110010100001000101010100;
		correct = 32'b10000010100010001001111110010110;
		#400; //1.2716532e-37 * -1.5786538 = -2.0075002e-37
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100011101000100100000101001;
		x2 = 32'b10100111001111010111011101010101;
		correct = 32'b11011100001101001100101100100101;
		#400; //7.7416017e+31 * -2.629371e-15 = -2.0355542e+17
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011011101111011110001110110010;
		x2 = 32'b11100010101100110100000011010110;
		correct = 32'b11111111000001001111011001001101;
		#400; //1.0689825e+17 * -1.6533196e+21 = -1.7673696e+38
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100111100001001001101100011000;
		x2 = 32'b00101100111001001101011110100001;
		correct = 32'b01010100111011010001001110100110;
		#400; //1.2524267e+24 * 6.5040894e-12 = 8145895000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000010111010110001111001111110;
		x2 = 32'b01000101110100110011111001110000;
		correct = 32'b10001001010000100000001101111010;
		#400; //-3.4547648e-37 * 6759.8047 = -2.3353535e-33
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111011101001110000000111000101;
		x2 = 32'b10101110100111111100011001110001;
		correct = 32'b10101010110100000111011100011101;
		#400; //0.0050966465 * -7.265733e-11 = -3.7030874e-13
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100010101100010011100101101111;
		x2 = 32'b10101100010011101001001101100011;
		correct = 32'b10001111100011110000001001000000;
		#400; //4.8036756e-18 * -2.9356177e-12 = -1.4101755e-29
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100001011101010111100001101;
		x2 = 32'b10001001111001100001110001101010;
		correct = 32'b00011110100111010000010010101001;
		#400; //-3001044700000.0 * -5.5397206e-33 = 1.6624949e-20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000111101100001010011010100111;
		x2 = 32'b00000110001011001011101001111010;
		correct = 32'b10001110011011100110000101001011;
		#400; //-90445.305 * 3.2486606e-35 = -2.938261e-30
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110111011100100010101110010111;
		x2 = 32'b11111011101111010011010001001010;
		correct = 32'b11110011101100101111101110100101;
		#400; //1.4434473e-05 * -1.9648093e+36 = -2.8360986e+31
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010011100101010101101011011010;
		x2 = 32'b00111110001011011000000010011101;
		correct = 32'b11010010010010100111001011011101;
		#400; //-1282948700000.0 * 0.16943593 = -217377620000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010000000000101011000010100010;
		x2 = 32'b00000000011010010100110001011000;
		correct = 32'b10010000110101110000010110101111;
		#400; //-8770456000.0 * 9.670114e-39 = -8.4811304e-29
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001001001100000111101000100;
		x2 = 32'b10100000000001100110111110101010;
		correct = 32'b00100001101011100110100011011001;
		#400; //-10.378727 * -1.1387188e-19 = 1.1818452e-18
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011000101011010010000011100011;
		x2 = 32'b11111110100011001001111100011111;
		correct = 32'b11010111101111100011001100110001;
		#400; //4.475266e-24 * -9.345906e+37 = -418254150000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100010000111011011000110001001;
		x2 = 32'b00110011011101111111001100001110;
		correct = 32'b10010110000110001011110000000011;
		#400; //-2.1371454e-18 * 5.7730226e-08 = -1.2337788e-25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110100100010101000111011000111;
		x2 = 32'b11000010100000000110101101010010;
		correct = 32'b11110111100010110000001011110011;
		#400; //8.782139e+31 * -64.20961 = -5.638977e+33
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100000011100010110111110100111;
		x2 = 32'b10100011000111000011011010110010;
		correct = 32'b10000100000100110101001110011111;
		#400; //2.0450437e-19 * -8.468359e-18 = -1.7318164e-36
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100110010100111111101010101011;
		x2 = 32'b00001101100100000111001111000101;
		correct = 32'b10110100011011110011100110111010;
		#400; //-2.5026083e+23 * 8.902556e-31 = -2.227961e-07
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110010000111111001100010010011;
		x2 = 32'b11101001110111100100011101011110;
		correct = 32'b01011100100010101001001011001101;
		#400; //-9.2897094e-09 * -3.358982e+25 = 3.1203965e+17
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100000100110011001111000001110;
		x2 = 32'b11001110100001111000001000101101;
		correct = 32'b00101111101000101010000011101101;
		#400; //-2.60238e-19 * -1136727700.0 = 2.9581973e-10
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111000100011101010100101011011;
		x2 = 32'b00000011001110111110111011111110;
		correct = 32'b00111100010100010111010111001001;
		#400; //2.314816e+34 * 5.522871e-37 = 0.01278443
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001000011010110110000000111;
		x2 = 32'b01110000101110000110101100001001;
		correct = 32'b11110010010010111100000110001100;
		#400; //-8.838874 * 4.565971e+29 = -4.0358042e+30
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101111001001010011100001110001;
		x2 = 32'b00010000011001111100101101110110;
		correct = 32'b11000000000101011001100100111110;
		#400; //-5.113326e+28 * 4.5713458e-29 = -2.3374782
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011101000100011001111010110010;
		x2 = 32'b00101100100100011001000010011101;
		correct = 32'b01001010001001011001101001001011;
		#400; //6.5581374e+17 * 4.137203e-12 = 2713234.8
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111001011110110001101110100011;
		x2 = 32'b01001010110000010000000110001111;
		correct = 32'b01000100101111010101000101011101;
		#400; //0.00023947521 * 6324423.5 = 1514.5426
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100111000001110001111111110010;
		x2 = 32'b00110000001011101000001001111100;
		correct = 32'b00010111101110000011100100101100;
		#400; //1.8752331e-15 * 6.348626e-10 = 1.1905154e-24
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010000010101011010011110010001;
		x2 = 32'b00010001001010011111111011101001;
		correct = 32'b10100010000011011110000001011101;
		#400; //-14338115000.0 * 1.34103e-28 = -1.922784e-18
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100110100011101001001111101;
		x2 = 32'b10111111100110100010101101111100;
		correct = 32'b01111100111111001011100010000110;
		#400; //-8.715674e+36 * -1.204452 = 1.0497611e+37
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110101000011001011000001101110;
		x2 = 32'b01110101101100110101010011110110;
		correct = 32'b11101011010001010001110000011100;
		#400; //-5.2410803e-07 * 4.5466033e+32 = -2.3829113e+26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000000100111001101110000101000;
		x2 = 32'b11100101010010011111100100110100;
		correct = 32'b11100110011101111000001100011011;
		#400; //4.9018745 * -5.961204e+22 = -2.9221075e+23
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110011100001000001111011101001;
		x2 = 32'b11010011011010010101001011001100;
		correct = 32'b11000111011100001101010110111011;
		#400; //6.1523515e-08 * -1002116500000.0 = -61653.73
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010011110010111101011110011111;
		x2 = 32'b00110001101101010111001110101010;
		correct = 32'b11000110000100000111101110001101;
		#400; //-1750991800000.0 * 5.280943e-09 = -9246.888
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110110111110011011011101011100;
		x2 = 32'b00011001111101100100110011011001;
		correct = 32'b11010001011100000100000100101001;
		#400; //-2.5324236e+33 * 2.5466842e-23 = -64492835000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01110011111010010101010010110011;
		x2 = 32'b00110111111001000111111101000000;
		correct = 32'b01101100010100000100001101101011;
		#400; //3.697275e+31 * 2.7238973e-05 = 1.0070998e+27
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101000011010010110010011010011;
		x2 = 32'b10001110000101000000100000100101;
		correct = 32'b10110111000001101111010110110111;
		#400; //4.408685e+24 * -1.824633e-30 = -8.044232e-06
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000101010101111000111100000010;
		x2 = 32'b01000101010011111111101101100001;
		correct = 32'b11001011001011110010000001001110;
		#400; //-3448.938 * 3327.7112 = -11477070.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011011011010000101000000001001;
		x2 = 32'b11101000111001110110111101110001;
		correct = 32'b01000100110100100000010101011001;
		#400; //-1.9216451e-22 * -8.743379e+24 = 1680.1671
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010110110010000110000010001010;
		x2 = 32'b00010101111100111110110101110100;
		correct = 32'b10101101001111101110110101111111;
		#400; //-110158480000000.0 * 9.8521553e-26 = -1.0852984e-11
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010000110110000011100011001010;
		x2 = 32'b01100011100001010101010100100001;
		correct = 32'b10110100111000010011101011001111;
		#400; //-8.5284475e-29 * 4.9191023e+21 = -4.1952305e-07
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111010101110011011100110010111;
		x2 = 32'b10001110110000010111101011010011;
		correct = 32'b01001010000011000101111000000110;
		#400; //-4.8216956e+35 * -4.769645e-30 = 2299777.5
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101011011011010100110110011011;
		x2 = 32'b01000100000001100011000101111111;
		correct = 32'b00101111111110001100100100000001;
		#400; //8.4307013e-13 * 536.7734 = 4.525376e-10
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011011011100100001100111110010;
		x2 = 32'b10000010110101000011011011111100;
		correct = 32'b10011110110010001011000101111100;
		#400; //6.814547e+16 * -3.118216e-37 = -2.124923e-20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01010000100100100111101010101010;
		x2 = 32'b01000101010011100001001100101011;
		correct = 32'b01010110011010111101001101011001;
		#400; //19660100000.0 * 3297.198 = 64823240000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110011100111011011000111101101;
		x2 = 32'b11000000101011111001001111100110;
		correct = 32'b10110100110110000100111101111000;
		#400; //7.343247e-08 * -5.486804 = -4.0290956e-07
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111100101010001000111010010101;
		x2 = 32'b01110100011111011001000110000000;
		correct = 32'b11110001101001101111010010110110;
		#400; //-0.0205758 * 8.035902e+31 = -1.6534512e+30
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001011100100011000100010011100;
		x2 = 32'b01001101011101100000101101111101;
		correct = 32'b01011001100010111101111111001110;
		#400; //19075384.0 * 257996750.0 = 4921387000000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001010011100000100001000101001;
		x2 = 32'b01001010001011001100000010011000;
		correct = 32'b01010101001000100010000100110100;
		#400; //3936394.2 * 2830374.0 = 11141468000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110100100100010111011110010100;
		x2 = 32'b00101101000010011010000101010010;
		correct = 32'b11100010000111000110100101010010;
		#400; //-9.220073e+31 * 7.823369e-12 = -7.213203e+20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110100101011011010111001001111;
		x2 = 32'b01101110011101101111111000001011;
		correct = 32'b01100011101001111001000111011010;
		#400; //3.2350587e-07 * 1.9110108e+28 = 6.182232e+21
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001110111100011000000011000010;
		x2 = 32'b00011111110100001101101111111011;
		correct = 32'b10101111010001010000100000100100;
		#400; //-2025873700.0 * 8.8455354e-20 = -1.7919938e-10
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000111110010100000100111100111;
		x2 = 32'b01001100110111011000111110011101;
		correct = 32'b11010101001011101101101111100100;
		#400; //-103443.805 * 116161770.0 = -12016215000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001010011000010000001011011001;
		x2 = 32'b01100010000111110010100100000001;
		correct = 32'b10101101000010111110010011001111;
		#400; //-1.08338915e-32 * 7.3399674e+20 = -7.952041e-12
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101110100000000111001111111010;
		x2 = 32'b00100010001000110100010011100100;
		correct = 32'b01010001001000111101100011010011;
		#400; //1.9877144e+28 * 2.212709e-18 = 43982336000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110011111110010111101110000001;
		x2 = 32'b10100011111011100101100000011110;
		correct = 32'b00011000011010000100011010110010;
		#400; //-1.1617431e-07 * -2.584133e-17 = 3.002099e-24
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101010111000111001011011001110;
		x2 = 32'b10001000100100010110011011101100;
		correct = 32'b00110100000000010100001111101011;
		#400; //-1.3756916e+26 * -8.751067e-34 = 1.203877e-07
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110011101011000110010011001100;
		x2 = 32'b00100110110101000001110011110010;
		correct = 32'b11011011000011101101011011110111;
		#400; //-2.7316878e+31 * 1.4718301e-15 = -4.0205803e+16
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11001011111011110010101110001110;
		x2 = 32'b11101110010001111101101101100001;
		correct = 32'b01111010101110101011011111010000;
		#400; //-31348508.0 * -1.5463182e+28 = 4.847477e+35
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011111001001101100101100011010;
		x2 = 32'b01011010111010100100000100011111;
		correct = 32'b10111010100110001010000000010100;
		#400; //-3.531987e-20 * 3.2968373e+16 = -0.0011644387
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110011000000110000001100001110;
		x2 = 32'b01101101111100100100110000001100;
		correct = 32'b11100001011101111111111110011101;
		#400; //-3.0503593e-08 * 9.3734134e+27 = -2.859228e+20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010100100110011110110000000000;
		x2 = 32'b11010010110101011101001001011010;
		correct = 32'b00101000000000001000111111010110;
		#400; //-1.5542138e-26 * -459178570000.0 = 7.136617e-15
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011111001000111110110111010101;
		x2 = 32'b00111110101001010110010011110011;
		correct = 32'b10011110010100111101000111011110;
		#400; //-3.4713323e-20 * 0.3230358 = -1.12136465e-20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011110010101000110110110110101;
		x2 = 32'b00100010111000100110010111010110;
		correct = 32'b01000001101110111101110101011011;
		#400; //3.8267724e+18 * 6.1365246e-18 = 23.483084
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001111101111100111001111101001;
		x2 = 32'b11001110100010111010000011111001;
		correct = 32'b00011110110011111100000101100010;
		#400; //-1.8780093e-29 * -1171291300.0 = 2.1996959e-20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011010001001110011000011011011;
		x2 = 32'b10100001010000111000011001010101;
		correct = 32'b10111011111111110110001111100100;
		#400; //1.176501e+16 * -6.6246357e-19 = -0.0077938903
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011010000110100000100101001;
		x2 = 32'b10000011011011110111101100101101;
		correct = 32'b00111111001101101010011111001000;
		#400; //-1.0138195e+36 * -7.0377186e-37 = 0.71349764
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000001000001101010101011111111;
		x2 = 32'b01000111011000001100100100101111;
		correct = 32'b10001000111011000111111011101000;
		#400; //-2.4734597e-38 * 57545.184 = -1.4233569e-33
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001010111100110100111110110110;
		x2 = 32'b00010100100101001111001001010111;
		correct = 32'b00100000000011011001000001101001;
		#400; //7972827.0 * 1.5039767e-26 = 1.1990946e-19
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101011110011101010010010110001;
		x2 = 32'b00111110111011101010010011010001;
		correct = 32'b11101011010000001010001000100111;
		#400; //-4.996329e+26 * 0.4661012 = -2.328795e+26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000000011100111011111011111;
		x2 = 32'b01000010101101011101100010110001;
		correct = 32'b10011011010010100110011010110001;
		#400; //-1.841359e-24 * 90.923225 = -1.674223e-22
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000100111111000000101011011101;
		x2 = 32'b01000100010100101001011001001011;
		correct = 32'b11001001110011110101010011100001;
		#400; //-2016.3395 * 842.3483 = -1698460.1
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01100001111011000110000001000000;
		x2 = 32'b10100000001000010011111010111110;
		correct = 32'b11000010100101001110001001110111;
		#400; //5.450459e+20 * -1.365799e-19 = -74.442314
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100000011000000001110000110011;
		x2 = 32'b00011111100010000010101010010000;
		correct = 32'b11000000011011100110100001111100;
		#400; //-6.4595354e+19 * 5.7668654e-20 = -3.7251272
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001011001000001101011100010101;
		x2 = 32'b01001000000101010111100000010110;
		correct = 32'b00010011101110111101000101000100;
		#400; //3.097669e-32 * 153056.34 = 4.741179e-27
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110001011101111001100100010000;
		x2 = 32'b10011101001110101010000010000100;
		correct = 32'b10001111001101001000000001110101;
		#400; //3.6030237e-09 * -2.469988e-21 = -8.899425e-30
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010100100001110101001111010001;
		x2 = 32'b11100011011110111011010000010111;
		correct = 32'b01111000100001010000111001100001;
		#400; //-4649814300000.0 * -4.6431096e+21 = 2.1589598e+34
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011010010101110010101111110101;
		x2 = 32'b11000001110100010100100111011111;
		correct = 32'b01011100101011111110100011111010;
		#400; //-1.5141363e+16 * -26.16107 = 3.9611425e+17
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101111111011101111110001011000;
		x2 = 32'b10001001110110100011101001001011;
		correct = 32'b10111010010010111011100101001110;
		#400; //1.4792499e+29 * -5.253641e-33 = -0.0007771448
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010000001110100111011001101001;
		x2 = 32'b11000011000111000001100100110010;
		correct = 32'b00010011111000110110010100000100;
		#400; //-3.6773252e-29 * -156.09842 = 5.7402465e-27
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10011000011101000001011011000001;
		x2 = 32'b01000000011111110000011111100100;
		correct = 32'b10011001011100110010101000110000;
		#400; //-3.1547749e-24 * 3.9848566 = -1.2571325e-23
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110001001010011001010010110001;
		x2 = 32'b11010010011100001100010000110010;
		correct = 32'b01000100000111110111110101011101;
		#400; //-2.4677258e-09 * -258520940000.0 = 637.9588
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010110101101000100101111111101;
		x2 = 32'b10100011011100110101011101001000;
		correct = 32'b00111010101010110110000110011010;
		#400; //-99119230000000.0 * -1.3191539e-17 = 0.0013075352
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001001111001010110100101111;
		x2 = 32'b10100111100000011101001011001110;
		correct = 32'b11100001001111110101110101000101;
		#400; //6.1229024e+34 * -3.6033247e-15 = -2.2062806e+20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11011111001011011101001110110101;
		x2 = 32'b01011000001101101100111010010101;
		correct = 32'b11110111111110000100000110010000;
		#400; //-1.2525554e+19 * 803993500000000.0 = -1.0070464e+34
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101111101011001100101110100110;
		x2 = 32'b10011010011011110010001111111101;
		correct = 32'b10001010101000010110101001101011;
		#400; //3.143132e-10 * -4.9453113e-23 = -1.5543766e-32
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11101000010001100000011001111001;
		x2 = 32'b00110100100101000001101111100100;
		correct = 32'b11011101011001010010001010100010;
		#400; //-3.7405919e+24 * 2.758744e-07 = -1.0319336e+18
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000001001101000001110111000001;
		x2 = 32'b10100110000111101100010010011001;
		correct = 32'b00100111110111110110100101011111;
		#400; //-11.257264 * -5.50837e-16 = 6.2009177e-15
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00001111011000010011010010001101;
		x2 = 32'b11001100001110000010000110110100;
		correct = 32'b10011100001000011111101101101011;
		#400; //1.11034774e-29 * -48269010.0 = -5.359538e-22
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111101111001011100001111111100;
		x2 = 32'b00110110011100111011100011111010;
		correct = 32'b00110100110110101011111100001101;
		#400; //0.11219022 * 3.6317492e-06 = 4.0744672e-07
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000000010110010011001011100111;
		x2 = 32'b10111110000010011010011110000100;
		correct = 32'b00111110111010011001010010111100;
		#400; //-3.3937318 * -0.13442808 = 0.45621288
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010010000101110100011000001010;
		x2 = 32'b11111011101000110000110001000100;
		correct = 32'b01001110010000001011000110110000;
		#400; //-4.773353e-28 * -1.6931863e+36 = 808217600.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100100010110000110101000111001;
		x2 = 32'b10100101000000011010110000000011;
		correct = 32'b00001001110110110011110111100001;
		#400; //-4.6927508e-17 * -1.1247246e-16 = 5.2780523e-33
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10010011101111100011010011110111;
		x2 = 32'b10111011110000000001010011100100;
		correct = 32'b00010000000011101011011100111111;
		#400; //-4.801497e-27 * -0.0058618654 = 2.814573e-29
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01101010010001111110100100100010;
		x2 = 32'b00110100010000101101010100110010;
		correct = 32'b01011111000110000010010100101000;
		#400; //6.0419294e+25 * 1.8145218e-07 = 1.0963213e+19
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011100011000011111011010101101;
		x2 = 32'b01010100011001001000000000010000;
		correct = 32'b01110001010010011011000010111100;
		#400; //2.5441237e+17 * 3925604300000.0 = 9.987223e+29
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10110000111101111011111000010010;
		x2 = 32'b10101010111011000110100011100000;
		correct = 32'b00011100011001001100100010110111;
		#400; //-1.8025637e-09 * -4.1994793e-13 = 7.569829e-22
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11010111001110000010101000011001;
		x2 = 32'b10101110010001101010001110010000;
		correct = 32'b01000110000011101110011000111010;
		#400; //-202490950000000.0 * -4.516526e-11 = 9145.557
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01011000101011011101100000100011;
		x2 = 32'b10110101111000001001011101101000;
		correct = 32'b11001111000110001000001111110000;
		#400; //1529150500000000.0 * -1.6733366e-06 = -2558783500.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111011110101110101011101100100;
		x2 = 32'b10101101110111101101001110110100;
		correct = 32'b01101010001110110110111111011101;
		#400; //-2.2362326e+36 * -2.5332493e-11 = 5.6649347e+25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000101100011010000101010111111;
		x2 = 32'b11010111010010000011110010110001;
		correct = 32'b11011101010111001010001110101011;
		#400; //4513.3433 * -220163000000000.0 = -9.936712e+17
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100011000000000101111001000001;
		x2 = 32'b11001111110000000110101011000010;
		correct = 32'b10110011010000001111100001110010;
		#400; //6.958853e-18 * -6456444000.0 = -4.4929443e-08
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001000111110010111000010111;
		x2 = 32'b00000110001110001101100101101101;
		correct = 32'b00111111111001011110000010100101;
		#400; //5.1656876e+34 * 3.4766293e-35 = 1.7959181
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000101100111010111010101100110;
		x2 = 32'b10011100111100001010101111100111;
		correct = 32'b00100011000101000000011111001011;
		#400; //-5038.675 * -1.5926303e-21 = 8.024746e-18
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010101011101000110011001001;
		x2 = 32'b00110111111000010111010101110110;
		correct = 32'b00111011000110011011100111010011;
		#400; //87.27497 * 2.6876787e-05 = 0.0023456707
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00010101101110100110110001110111;
		x2 = 32'b01100111101111101110110100111001;
		correct = 32'b00111110000010110000100101000000;
		#400; //7.529593e-26 * 1.8032512e+24 = 0.13577747
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000110000101110001101001110001;
		x2 = 32'b00010100100100101110111111011010;
		correct = 32'b00011011001011010111010101001110;
		#400; //9670.61 * 1.4836837e-26 = 1.4348128e-22
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00000100101100111000101000110001;
		x2 = 32'b01010010001100011111100011001100;
		correct = 32'b00010111011110011010001000010010;
		#400; //4.2209607e-36 * 191095830000.0 = 8.06608e-25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11100001000010001001001000011010;
		x2 = 32'b10010001011011000011001010001000;
		correct = 32'b00110010111111000000001101001010;
		#400; //-1.574553e+20 * -1.8632689e-28 = 2.9338157e-08
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100100110011000101010100111100;
		x2 = 32'b01011100110000010011111010000000;
		correct = 32'b01000010000110100011111000100101;
		#400; //8.861529e-17 * 4.3514712e+17 = 38.560688
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100101101110000001101000101111;
		x2 = 32'b11010111000000101010110101010110;
		correct = 32'b00111101001110111111001111100111;
		#400; //-3.1936655e-16 * -143680980000000.0 = 0.0458869
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000100011000001100001100011101;
		x2 = 32'b00101101000011001010110110000001;
		correct = 32'b00110001111101110000011000010010;
		#400; //899.04865 * 7.996604e-12 = 7.1893362e-09
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11110111010000101000000110110111;
		x2 = 32'b00001010000010110100001111100011;
		correct = 32'b11000001110100111010000000000110;
		#400; //-3.9450645e+33 * 6.7053746e-33 = -26.453136
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00100101000000010001100010000101;
		x2 = 32'b11100100110111101011110001000000;
		correct = 32'b11001010011000001010010001100011;
		#400; //1.1197274e-16 * -3.2869936e+22 = -3680536.8
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10001110110010011010111010011000;
		x2 = 32'b11001011011101011110101010010010;
		correct = 32'b00011010110000011011110011100100;
		#400; //-4.9718453e-30 * -16116370.0 = 8.01281e-23
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10100000001111011010010000001001;
		x2 = 32'b01110001000111011001101011011101;
		correct = 32'b11010001111010011000000010100100;
		#400; //-1.6063197e-19 * 7.804218e+29 = -125360700000.0
					end  
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111100100011111001001111010010;
		x2 = 32'b00001100100011000011010110011110;
		correct = 32'b00001001100111010100010111010010;
		#400; //0.01752654 * 2.1602685e-31 = 3.7862034e-33
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10000011001010101000100001100011;
		x2 = 32'b11011111001101100111000001010001;
		correct = 32'b00100010111100110000111110010000;
		#400; //-5.0115074e-37 * -1.3146096e+19 = 6.588176e-18
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000010111101111110010110011101;
		x2 = 32'b01011101100010001111101010101001;
		correct = 32'b01100001000001001010010010110101;
		#400; //123.94846 * 1.2337984e+18 = 1.5292741e+20
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11111100001010001010111101100001;
		x2 = 32'b10111101100010010101110111010010;
		correct = 32'b01111010001101010000011101011010;
		#400; //-3.503452e+36 * -0.06707348 = 2.349887e+35
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111011001000110001001010111011;
		x2 = 32'b10101100101011000001101110111100;
		correct = 32'b11101000010110110100010010000001;
		#400; //8.467243e+35 * -4.891613e-12 = -4.1418477e+24
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10111110101011111101001101001110;
		x2 = 32'b11101011000011001110100001100111;
		correct = 32'b01101010010000011000111001011010;
		#400; //-0.343409 * -1.703471e+26 = 5.849873e+25
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b10101001000100110100111001001100;
		x2 = 32'b01000101011100011110111001111111;
		correct = 32'b10101111000010110011010111110001;
		#400; //-3.270847e-14 * 3870.906 = -1.266114e-10
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00110101010100111000010101010000;
		x2 = 32'b00111101010100011010010010010001;
		correct = 32'b00110011001011010011011111010000;
		#400; //7.879762e-07 * 0.051182333 = 4.0330463e-08
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01000000111011000010000100000111;
		x2 = 32'b10001010010000101110010010100111;
		correct = 32'b10001011101100111100001111101111;
		#400; //7.3790317 * -9.383765e-33 = -6.92431e-32
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00011000010110010100010001000110;
		x2 = 32'b11011011100010110011011011000110;
		correct = 32'b10110100011011000100110100011101;
		#400; //2.8081062e-24 * -7.837049e+16 = -2.2007266e-07
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001010110100110000110011111011;
		x2 = 32'b11011100000001100011100000011010;
		correct = 32'b11100111010111010100111000010111;
		#400; //6915709.5 * -1.5111732e+17 = -1.0450835e+24
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b11000011100110011111110100111100;
		x2 = 32'b10010001000111101111101011100001;
		correct = 32'b00010101001111110100001001100111;
		#400; //-307.9784 * -1.254131e-28 = 3.8624525e-26
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00101001110001010111101110101010;
		x2 = 32'b11000111111000100011000010001110;
		correct = 32'b10110010001011100111110010100001;
		#400; //8.77001e-14 * -115809.11 = -1.015647e-08
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01001100001010111011011011011101;
		x2 = 32'b11000010011001101101010001110111;
		correct = 32'b11001111000110101101010011001110;
		#400; //45013876.0 * -57.707485 = -2597637600.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b01111001010011001100011000011001;
		x2 = 32'b10000000110110001110101111100100;
		correct = 32'b10111010101011011000001111010101;
		#400; //6.6452904e+34 * -1.9921089e-38 = -0.0013238142
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		x1 = 32'b00111110111111110100010010100101;
		x2 = 32'b01010110101110100001000101111001;
		correct = 32'b01010110001110011000100101001100;
		#400; //0.4985706 * 102292100000000.0 = 50999834000000.0
					end 
 begin
			$display ("A      : %x2 %x2 %x2", x1[31], x1[30:23], x1[22:0]);
			$display ("B      : %x2 %x2 %x2", x2[31], x2[30:23], x2[22:0]);
			$display ("Output : %x2 %x2 %x2", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end
end
endmodule